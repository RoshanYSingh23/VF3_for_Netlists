module c1355(inout G1, inout G10, inout G11, inout G12, inout G13, inout N384, inout N385, inout N386, inout N387, inout N388, inout N389, inout N390, inout N391, inout N392, inout N393, inout N394, inout N395, inout N396, inout N397, inout N398, inout N399, inout N400, inout N401, inout N402, inout N403, inout N404, inout N405, inout N406, inout N407, inout N408, inout N409, inout N410, inout N411, inout N412, inout N413, inout N414, inout N415, inout G14, inout G15, inout G16, inout G17, inout G18, inout G19, inout G2, inout G20, inout G21, inout G22, inout G23, inout G24, inout G25, inout G26, inout G27, inout G28, inout G29, inout G3, inout G30, inout G31, inout G32, inout G33, inout G34, inout G35, inout G36, inout G37, inout G38, inout G39, inout G4, inout G40, inout G41, inout G5, inout G6, inout G7, inout G8, inout G9, inout VDD, inout GND)
	INVX1 X1 (.VDD(VDD), .GND(), .A(n230), .Y(U254/a_2_6#));
	INVX1 X2 (.VDD(), .GND(), .A(n232), .Y());
	INVX1 X3 (.VDD(VDD), .GND(GND), .A(U254/a_2_6#), .Y(n305));
	INVX1 X4 (.VDD(VDD), .GND(), .A(n231), .Y(U255/a_2_6#));
	INVX1 X5 (.VDD(), .GND(), .A(n233), .Y());
	INVX1 X6 (.VDD(VDD), .GND(GND), .A(U255/a_2_6#), .Y(n350));
	INVX1 X7 (.VDD(), .GND(), .A(n293), .Y());
	INVX1 X8 (.VDD(VDD), .GND(GND), .A(U256/a_2_6#), .Y(n222));
	INVX1 X9 (.VDD(), .GND(), .A(n304), .Y());
	INVX1 X10 (.VDD(VDD), .GND(GND), .A(U257/a_2_6#), .Y(n223));
	INVX1 X11 (.VDD(), .GND(), .A(n314), .Y());
	INVX1 X12 (.VDD(VDD), .GND(GND), .A(U258/a_2_6#), .Y(n224));
	INVX1 X13 (.VDD(), .GND(), .A(n323), .Y());
	INVX1 X14 (.VDD(VDD), .GND(GND), .A(U259/a_2_6#), .Y(n225));
	INVX1 X15 (.VDD(), .GND(), .A(n341), .Y());
	INVX1 X16 (.VDD(VDD), .GND(GND), .A(U260/a_2_6#), .Y(n226));
	INVX1 X17 (.VDD(), .GND(), .A(n349), .Y());
	INVX1 X18 (.VDD(VDD), .GND(GND), .A(U261/a_2_6#), .Y(n227));
	INVX1 X19 (.VDD(), .GND(), .A(n358), .Y());
	INVX1 X20 (.VDD(VDD), .GND(GND), .A(U262/a_2_6#), .Y(n228));
	INVX1 X21 (.VDD(), .GND(), .A(n365), .Y());
	INVX1 X22 (.VDD(VDD), .GND(GND), .A(U263/a_2_6#), .Y(n229));
	INVX1 X23 (.VDD(), .GND(), .A(n325), .Y());
	INVX1 X24 (.VDD(VDD), .GND(GND), .A(U264/a_2_6#), .Y(n230));
	INVX1 X25 (.VDD(), .GND(), .A(n375), .Y());
	INVX1 X26 (.VDD(VDD), .GND(GND), .A(U265/a_2_6#), .Y(n231));
	INVX1 X27 (.VDD(), .GND(), .A(n326), .Y());
	INVX1 X28 (.VDD(VDD), .GND(GND), .A(U266/a_2_6#), .Y(n232));
	INVX1 X29 (.VDD(), .GND(), .A(n376), .Y());
	INVX1 X30 (.VDD(VDD), .GND(GND), .A(U267/a_2_6#), .Y(n233));
	INVX1 X31 (.VDD(), .GND(GND), .A(n307), .Y(U268/a_2_54#));
	INVX1 X32 (.VDD(), .GND(), .A(n276), .Y());
	INVX1 X33 (.VDD(VDD), .GND(GND), .A(U268/a_2_54#), .Y(n306));
	INVX1 X34 (.VDD(VDD), .GND(GND), .A(n306), .Y(n234));
	INVX1 X35 (.VDD(), .GND(GND), .A(n316), .Y(U270/a_2_54#));
	INVX1 X36 (.VDD(), .GND(), .A(n282), .Y());
	INVX1 X37 (.VDD(VDD), .GND(GND), .A(U270/a_2_54#), .Y(n315));
	INVX1 X38 (.VDD(VDD), .GND(GND), .A(n315), .Y(n235));
	INVX1 X39 (.VDD(), .GND(GND), .A(n286), .Y(U272/a_2_54#));
	INVX1 X40 (.VDD(), .GND(), .A(n277), .Y());
	INVX1 X41 (.VDD(VDD), .GND(GND), .A(U272/a_2_54#), .Y(n351));
	INVX1 X42 (.VDD(VDD), .GND(GND), .A(n351), .Y(n236));
	INVX1 X43 (.VDD(), .GND(GND), .A(n288), .Y(U274/a_2_54#));
	INVX1 X44 (.VDD(), .GND(), .A(n283), .Y());
	INVX1 X45 (.VDD(VDD), .GND(GND), .A(U274/a_2_54#), .Y(n359));
	INVX1 X46 (.VDD(VDD), .GND(GND), .A(n359), .Y(n237));
	INVX1 X47 (.VDD(VDD), .GND(GND), .A(n305), .Y(n238));
	INVX1 X48 (.VDD(VDD), .GND(GND), .A(n350), .Y(n239));
	INVX1 X49 (.VDD(VDD), .GND(), .A(n353), .Y(U278/a_2_6#));
	INVX1 X50 (.VDD(), .GND(), .A(n340), .Y());
	INVX1 X51 (.VDD(VDD), .GND(GND), .A(U278/a_2_6#), .Y(n356));
	INVX1 X52 (.VDD(VDD), .GND(GND), .A(n356), .Y(n240));
	INVX1 X53 (.VDD(VDD), .GND(), .A(n344), .Y(U280/a_2_6#));
	INVX1 X54 (.VDD(), .GND(), .A(n316), .Y());
	INVX1 X55 (.VDD(VDD), .GND(GND), .A(U280/a_2_6#), .Y(n346));
	INVX1 X56 (.VDD(VDD), .GND(GND), .A(n346), .Y(n241));
	INVX1 X57 (.VDD(VDD), .GND(), .A(G36), .Y(U282/a_2_6#));
	INVX1 X58 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X59 (.VDD(VDD), .GND(GND), .A(U282/a_2_6#), .Y(n391));
	INVX1 X60 (.VDD(VDD), .GND(GND), .A(n391), .Y(n242));
	INVX1 X61 (.VDD(VDD), .GND(), .A(G38), .Y(U284/a_2_6#));
	INVX1 X62 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X63 (.VDD(VDD), .GND(GND), .A(U284/a_2_6#), .Y(n438));
	INVX1 X64 (.VDD(VDD), .GND(GND), .A(n438), .Y(n243));
	INVX1 X65 (.VDD(VDD), .GND(), .A(G37), .Y(U286/a_2_6#));
	INVX1 X66 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X67 (.VDD(VDD), .GND(GND), .A(U286/a_2_6#), .Y(n420));
	INVX1 X68 (.VDD(VDD), .GND(GND), .A(n420), .Y(n244));
	INVX1 X69 (.VDD(VDD), .GND(), .A(G40), .Y(U288/a_2_6#));
	INVX1 X70 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X71 (.VDD(VDD), .GND(GND), .A(U288/a_2_6#), .Y(n429));
	INVX1 X72 (.VDD(VDD), .GND(GND), .A(n429), .Y(n245));
	INVX1 X73 (.VDD(VDD), .GND(), .A(n361), .Y(U290/a_2_6#));
	INVX1 X74 (.VDD(), .GND(), .A(n336), .Y());
	INVX1 X75 (.VDD(VDD), .GND(GND), .A(U290/a_2_6#), .Y(n362));
	INVX1 X76 (.VDD(VDD), .GND(GND), .A(n362), .Y(n246));
	INVX1 X77 (.VDD(VDD), .GND(), .A(n319), .Y(U292/a_2_6#));
	INVX1 X78 (.VDD(), .GND(), .A(n288), .Y());
	INVX1 X79 (.VDD(VDD), .GND(GND), .A(U292/a_2_6#), .Y(n320));
	INVX1 X80 (.VDD(VDD), .GND(GND), .A(n320), .Y(n247));
	INVX1 X81 (.VDD(VDD), .GND(), .A(G41), .Y(U294/a_2_6#));
	INVX1 X82 (.VDD(), .GND(), .A(G39), .Y());
	INVX1 X83 (.VDD(VDD), .GND(GND), .A(U294/a_2_6#), .Y(n373));
	INVX1 X84 (.VDD(VDD), .GND(GND), .A(n373), .Y(n248));
	INVX1 X85 (.VDD(VDD), .GND(), .A(G35), .Y(U296/a_2_6#));
	INVX1 X86 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X87 (.VDD(VDD), .GND(GND), .A(U296/a_2_6#), .Y(n410));
	INVX1 X88 (.VDD(VDD), .GND(GND), .A(n410), .Y(n249));
	INVX1 X89 (.VDD(VDD), .GND(), .A(n361), .Y(U298/a_2_6#));
	INVX1 X90 (.VDD(), .GND(), .A(n307), .Y());
	INVX1 X91 (.VDD(VDD), .GND(GND), .A(U298/a_2_6#), .Y(n360));
	INVX1 X92 (.VDD(VDD), .GND(GND), .A(n360), .Y(n250));
	INVX1 X93 (.VDD(VDD), .GND(), .A(n353), .Y(U300/a_2_6#));
	INVX1 X94 (.VDD(), .GND(), .A(n316), .Y());
	INVX1 X95 (.VDD(VDD), .GND(GND), .A(U300/a_2_6#), .Y(n355));
	INVX1 X96 (.VDD(VDD), .GND(GND), .A(n355), .Y(n251));
	INVX1 X97 (.VDD(VDD), .GND(), .A(n344), .Y(U302/a_2_6#));
	INVX1 X98 (.VDD(), .GND(), .A(n340), .Y());
	INVX1 X99 (.VDD(VDD), .GND(GND), .A(U302/a_2_6#), .Y(n348));
	INVX1 X100 (.VDD(VDD), .GND(GND), .A(n348), .Y(n252));
	INVX1 X101 (.VDD(VDD), .GND(), .A(n319), .Y(U304/a_2_6#));
	INVX1 X102 (.VDD(), .GND(), .A(n286), .Y());
	INVX1 X103 (.VDD(VDD), .GND(GND), .A(U304/a_2_6#), .Y(n318));
	INVX1 X104 (.VDD(VDD), .GND(GND), .A(n318), .Y(n253));
	INVX1 X105 (.VDD(VDD), .GND(), .A(n310), .Y(U306/a_2_6#));
	INVX1 X106 (.VDD(), .GND(), .A(n290), .Y());
	INVX1 X107 (.VDD(VDD), .GND(GND), .A(U306/a_2_6#), .Y(n312));
	INVX1 X108 (.VDD(VDD), .GND(GND), .A(n312), .Y(n254));
	INVX1 X109 (.VDD(VDD), .GND(), .A(n300), .Y(U308/a_2_6#));
	INVX1 X110 (.VDD(), .GND(), .A(n292), .Y());
	INVX1 X111 (.VDD(VDD), .GND(GND), .A(U308/a_2_6#), .Y(n303));
	INVX1 X112 (.VDD(VDD), .GND(GND), .A(n303), .Y(n255));
	INVX1 X113 (.VDD(VDD), .GND(), .A(n334), .Y(U310/a_2_6#));
	INVX1 X114 (.VDD(), .GND(), .A(n340), .Y());
	INVX1 X115 (.VDD(VDD), .GND(GND), .A(U310/a_2_6#), .Y(n338));
	INVX1 X116 (.VDD(VDD), .GND(GND), .A(n338), .Y(n256));
	INVX1 X117 (.VDD(VDD), .GND(), .A(G34), .Y(U312/a_2_6#));
	INVX1 X118 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X119 (.VDD(VDD), .GND(GND), .A(U312/a_2_6#), .Y(n383));
	INVX1 X120 (.VDD(VDD), .GND(GND), .A(n383), .Y(n257));
	INVX1 X121 (.VDD(VDD), .GND(), .A(n353), .Y(U314/a_2_6#));
	INVX1 X122 (.VDD(), .GND(), .A(n307), .Y());
	INVX1 X123 (.VDD(VDD), .GND(GND), .A(U314/a_2_6#), .Y(n352));
	INVX1 X124 (.VDD(VDD), .GND(GND), .A(n352), .Y(n258));
	INVX1 X125 (.VDD(VDD), .GND(), .A(n344), .Y(U316/a_2_6#));
	INVX1 X126 (.VDD(), .GND(), .A(n336), .Y());
	INVX1 X127 (.VDD(VDD), .GND(GND), .A(U316/a_2_6#), .Y(n345));
	INVX1 X128 (.VDD(VDD), .GND(GND), .A(n345), .Y(n259));
	INVX1 X129 (.VDD(VDD), .GND(), .A(n319), .Y(U318/a_2_6#));
	INVX1 X130 (.VDD(), .GND(), .A(n290), .Y());
	INVX1 X131 (.VDD(VDD), .GND(GND), .A(U318/a_2_6#), .Y(n321));
	INVX1 X132 (.VDD(VDD), .GND(GND), .A(n321), .Y(n260));
	INVX1 X133 (.VDD(VDD), .GND(), .A(n310), .Y(U320/a_2_6#));
	INVX1 X134 (.VDD(), .GND(), .A(n286), .Y());
	INVX1 X135 (.VDD(VDD), .GND(GND), .A(U320/a_2_6#), .Y(n309));
	INVX1 X136 (.VDD(VDD), .GND(GND), .A(n309), .Y(n261));
	INVX1 X137 (.VDD(VDD), .GND(), .A(n300), .Y(U322/a_2_6#));
	INVX1 X138 (.VDD(), .GND(), .A(n288), .Y());
	INVX1 X139 (.VDD(VDD), .GND(GND), .A(U322/a_2_6#), .Y(n301));
	INVX1 X140 (.VDD(VDD), .GND(GND), .A(n301), .Y(n262));
	INVX1 X141 (.VDD(VDD), .GND(), .A(n285), .Y(U324/a_2_6#));
	INVX1 X142 (.VDD(), .GND(), .A(n292), .Y());
	INVX1 X143 (.VDD(VDD), .GND(GND), .A(U324/a_2_6#), .Y(n291));
	INVX1 X144 (.VDD(VDD), .GND(GND), .A(n291), .Y(n263));
	INVX1 X145 (.VDD(VDD), .GND(), .A(G33), .Y(U326/a_2_6#));
	INVX1 X146 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X147 (.VDD(VDD), .GND(GND), .A(U326/a_2_6#), .Y(n400));
	INVX1 X148 (.VDD(VDD), .GND(GND), .A(n400), .Y(n264));
	INVX1 X149 (.VDD(VDD), .GND(), .A(n353), .Y(U328/a_2_6#));
	INVX1 X150 (.VDD(), .GND(), .A(n336), .Y());
	INVX1 X151 (.VDD(VDD), .GND(GND), .A(U328/a_2_6#), .Y(n354));
	INVX1 X152 (.VDD(VDD), .GND(GND), .A(n354), .Y(n265));
	INVX1 X153 (.VDD(VDD), .GND(), .A(n344), .Y(U330/a_2_6#));
	INVX1 X154 (.VDD(), .GND(), .A(n307), .Y());
	INVX1 X155 (.VDD(VDD), .GND(GND), .A(U330/a_2_6#), .Y(n343));
	INVX1 X156 (.VDD(VDD), .GND(GND), .A(n343), .Y(n266));
	INVX1 X157 (.VDD(VDD), .GND(), .A(n334), .Y(U332/a_2_6#));
	INVX1 X158 (.VDD(), .GND(), .A(n316), .Y());
	INVX1 X159 (.VDD(VDD), .GND(GND), .A(U332/a_2_6#), .Y(n337));
	INVX1 X160 (.VDD(VDD), .GND(GND), .A(n337), .Y(n267));
	INVX1 X161 (.VDD(VDD), .GND(), .A(n319), .Y(U334/a_2_6#));
	INVX1 X162 (.VDD(), .GND(), .A(n292), .Y());
	INVX1 X163 (.VDD(VDD), .GND(GND), .A(U334/a_2_6#), .Y(n322));
	INVX1 X164 (.VDD(VDD), .GND(GND), .A(n322), .Y(n268));
	INVX1 X165 (.VDD(VDD), .GND(), .A(n310), .Y(U336/a_2_6#));
	INVX1 X166 (.VDD(), .GND(), .A(n288), .Y());
	INVX1 X167 (.VDD(VDD), .GND(GND), .A(U336/a_2_6#), .Y(n311));
	INVX1 X168 (.VDD(VDD), .GND(GND), .A(n311), .Y(n269));
	INVX1 X169 (.VDD(VDD), .GND(), .A(n300), .Y(U338/a_2_6#));
	INVX1 X170 (.VDD(), .GND(), .A(n286), .Y());
	INVX1 X171 (.VDD(VDD), .GND(GND), .A(U338/a_2_6#), .Y(n299));
	INVX1 X172 (.VDD(VDD), .GND(GND), .A(n299), .Y(n270));
	INVX1 X173 (.VDD(VDD), .GND(), .A(n285), .Y(U340/a_2_6#));
	INVX1 X174 (.VDD(), .GND(), .A(n290), .Y());
	INVX1 X175 (.VDD(VDD), .GND(GND), .A(U340/a_2_6#), .Y(n289));
	INVX1 X176 (.VDD(VDD), .GND(GND), .A(n289), .Y(n271));
	INVX1 X177 (.VDD(VDD), .GND(), .A(n361), .Y(U342/a_2_6#));
	INVX1 X178 (.VDD(), .GND(), .A(n340), .Y());
	INVX1 X179 (.VDD(VDD), .GND(GND), .A(U342/a_2_6#), .Y(n364));
	INVX1 X180 (.VDD(VDD), .GND(GND), .A(n364), .Y(n272));
	INVX1 X181 (.VDD(VDD), .GND(), .A(n334), .Y(U344/a_2_6#));
	INVX1 X182 (.VDD(), .GND(), .A(n307), .Y());
	INVX1 X183 (.VDD(VDD), .GND(GND), .A(U344/a_2_6#), .Y(n333));
	INVX1 X184 (.VDD(VDD), .GND(GND), .A(n333), .Y(n273));
	INVX1 X185 (.VDD(VDD), .GND(), .A(n310), .Y(U346/a_2_6#));
	INVX1 X186 (.VDD(), .GND(), .A(n292), .Y());
	INVX1 X187 (.VDD(VDD), .GND(GND), .A(U346/a_2_6#), .Y(n313));
	INVX1 X188 (.VDD(VDD), .GND(GND), .A(n313), .Y(n274));
	INVX1 X189 (.VDD(VDD), .GND(), .A(n285), .Y(U348/a_2_6#));
	INVX1 X190 (.VDD(), .GND(), .A(n286), .Y());
	INVX1 X191 (.VDD(VDD), .GND(GND), .A(U348/a_2_6#), .Y(n284));
	INVX1 X192 (.VDD(VDD), .GND(GND), .A(n284), .Y(n275));
	INVX1 X193 (.VDD(VDD), .GND(), .A(n336), .Y(U350/a_2_6#));
	INVX1 X194 (.VDD(), .GND(), .A(n316), .Y());
	INVX1 X195 (.VDD(VDD), .GND(GND), .A(U350/a_2_6#), .Y(n308));
	INVX1 X196 (.VDD(VDD), .GND(GND), .A(n308), .Y(n276));
	INVX1 X197 (.VDD(VDD), .GND(), .A(n290), .Y(U352/a_2_6#));
	INVX1 X198 (.VDD(), .GND(), .A(n288), .Y());
	INVX1 X199 (.VDD(VDD), .GND(GND), .A(U352/a_2_6#), .Y(n328));
	INVX1 X200 (.VDD(VDD), .GND(GND), .A(n328), .Y(n277));
	INVX1 X201 (.VDD(VDD), .GND(), .A(n361), .Y(U354/a_2_6#));
	INVX1 X202 (.VDD(), .GND(), .A(n316), .Y());
	INVX1 X203 (.VDD(VDD), .GND(GND), .A(U354/a_2_6#), .Y(n363));
	INVX1 X204 (.VDD(VDD), .GND(GND), .A(n363), .Y(n278));
	INVX1 X205 (.VDD(VDD), .GND(), .A(n334), .Y(U356/a_2_6#));
	INVX1 X206 (.VDD(), .GND(), .A(n336), .Y());
	INVX1 X207 (.VDD(VDD), .GND(GND), .A(U356/a_2_6#), .Y(n335));
	INVX1 X208 (.VDD(VDD), .GND(GND), .A(n335), .Y(n279));
	INVX1 X209 (.VDD(VDD), .GND(), .A(n300), .Y(U358/a_2_6#));
	INVX1 X210 (.VDD(), .GND(), .A(n290), .Y());
	INVX1 X211 (.VDD(VDD), .GND(GND), .A(U358/a_2_6#), .Y(n302));
	INVX1 X212 (.VDD(VDD), .GND(GND), .A(n302), .Y(n280));
	INVX1 X213 (.VDD(VDD), .GND(), .A(n285), .Y(U360/a_2_6#));
	INVX1 X214 (.VDD(), .GND(), .A(n288), .Y());
	INVX1 X215 (.VDD(VDD), .GND(GND), .A(U360/a_2_6#), .Y(n287));
	INVX1 X216 (.VDD(VDD), .GND(GND), .A(n287), .Y(n281));
	INVX1 X217 (.VDD(VDD), .GND(), .A(n340), .Y(U362/a_2_6#));
	INVX1 X218 (.VDD(), .GND(), .A(n307), .Y());
	INVX1 X219 (.VDD(VDD), .GND(GND), .A(U362/a_2_6#), .Y(n317));
	INVX1 X220 (.VDD(VDD), .GND(GND), .A(n317), .Y(n282));
	INVX1 X221 (.VDD(VDD), .GND(), .A(n292), .Y(U364/a_2_6#));
	INVX1 X222 (.VDD(), .GND(), .A(n286), .Y());
	INVX1 X223 (.VDD(VDD), .GND(GND), .A(U364/a_2_6#), .Y(n331));
	INVX1 X224 (.VDD(VDD), .GND(GND), .A(n331), .Y(n283));
	INVX1 X225 (.VDD(), .GND(), .A(n275), .Y());
	INVX1 X226 (.VDD(VDD), .GND(GND), .A(U366/a_13_43#), .Y(U366/a_18_54#));
	INVX1 X227 (.VDD(), .GND(), .A(n275), .Y());
	INVX1 X228 (.VDD(), .GND(), .A(U366/a_2_6#), .Y());
	INVX1 X229 (.VDD(), .GND(), .A(G32), .Y());
	INVX1 X230 (.VDD(VDD), .GND(GND), .A(G32), .Y(U366/a_13_43#));
	INVX1 X231 (.VDD(), .GND(), .A(n281), .Y());
	INVX1 X232 (.VDD(VDD), .GND(GND), .A(U367/a_13_43#), .Y(U367/a_18_54#));
	INVX1 X233 (.VDD(), .GND(), .A(n281), .Y());
	INVX1 X234 (.VDD(), .GND(), .A(U367/a_2_6#), .Y());
	INVX1 X235 (.VDD(), .GND(), .A(G31), .Y());
	INVX1 X236 (.VDD(VDD), .GND(GND), .A(G31), .Y(U367/a_13_43#));
	INVX1 X237 (.VDD(), .GND(), .A(n271), .Y());
	INVX1 X238 (.VDD(VDD), .GND(GND), .A(U368/a_13_43#), .Y(U368/a_18_54#));
	INVX1 X239 (.VDD(), .GND(), .A(n271), .Y());
	INVX1 X240 (.VDD(), .GND(), .A(U368/a_2_6#), .Y());
	INVX1 X241 (.VDD(), .GND(), .A(G30), .Y());
	INVX1 X242 (.VDD(VDD), .GND(GND), .A(G30), .Y(U368/a_13_43#));
	INVX1 X243 (.VDD(), .GND(), .A(n263), .Y());
	INVX1 X244 (.VDD(VDD), .GND(GND), .A(U369/a_13_43#), .Y(U369/a_18_54#));
	INVX1 X245 (.VDD(), .GND(), .A(n263), .Y());
	INVX1 X246 (.VDD(), .GND(), .A(U369/a_2_6#), .Y());
	INVX1 X247 (.VDD(), .GND(), .A(G29), .Y());
	INVX1 X248 (.VDD(VDD), .GND(GND), .A(G29), .Y(U369/a_13_43#));
	INVX1 X249 (.VDD(VDD), .GND(GND), .A(n222), .Y(n285));
	INVX1 X250 (.VDD(VDD), .GND(GND), .A(n294), .Y(n293));
	INVX1 X251 (.VDD(), .GND(), .A(n295), .Y());
	INVX1 X252 (.VDD(VDD), .GND(), .A(n296), .Y(n293));
	INVX1 X253 (.VDD(), .GND(GND), .A(n297), .Y(n296));
	INVX1 X254 (.VDD(VDD), .GND(GND), .A(n297), .Y(U372/a_2_64#));
	INVX1 X255 (.VDD(), .GND(), .A(n305), .Y());
	INVX1 X256 (.VDD(), .GND(), .A(n305), .Y());
	INVX1 X257 (.VDD(), .GND(GND), .A(n298), .Y(n296));
	INVX1 X258 (.VDD(), .GND(), .A(n298), .Y());
	INVX1 X259 (.VDD(), .GND(), .A(n270), .Y());
	INVX1 X260 (.VDD(VDD), .GND(GND), .A(U373/a_13_43#), .Y(U373/a_18_54#));
	INVX1 X261 (.VDD(), .GND(), .A(n270), .Y());
	INVX1 X262 (.VDD(), .GND(), .A(U373/a_2_6#), .Y());
	INVX1 X263 (.VDD(), .GND(), .A(G28), .Y());
	INVX1 X264 (.VDD(VDD), .GND(GND), .A(G28), .Y(U373/a_13_43#));
	INVX1 X265 (.VDD(), .GND(), .A(n262), .Y());
	INVX1 X266 (.VDD(VDD), .GND(GND), .A(U374/a_13_43#), .Y(U374/a_18_54#));
	INVX1 X267 (.VDD(), .GND(), .A(n262), .Y());
	INVX1 X268 (.VDD(), .GND(), .A(U374/a_2_6#), .Y());
	INVX1 X269 (.VDD(), .GND(), .A(G27), .Y());
	INVX1 X270 (.VDD(VDD), .GND(GND), .A(G27), .Y(U374/a_13_43#));
	INVX1 X271 (.VDD(), .GND(), .A(n280), .Y());
	INVX1 X272 (.VDD(VDD), .GND(GND), .A(U375/a_13_43#), .Y(U375/a_18_54#));
	INVX1 X273 (.VDD(), .GND(), .A(n280), .Y());
	INVX1 X274 (.VDD(), .GND(), .A(U375/a_2_6#), .Y());
	INVX1 X275 (.VDD(), .GND(), .A(G26), .Y());
	INVX1 X276 (.VDD(VDD), .GND(GND), .A(G26), .Y(U375/a_13_43#));
	INVX1 X277 (.VDD(), .GND(), .A(n255), .Y());
	INVX1 X278 (.VDD(VDD), .GND(GND), .A(U376/a_13_43#), .Y(U376/a_18_54#));
	INVX1 X279 (.VDD(), .GND(), .A(n255), .Y());
	INVX1 X280 (.VDD(), .GND(), .A(U376/a_2_6#), .Y());
	INVX1 X281 (.VDD(), .GND(), .A(G25), .Y());
	INVX1 X282 (.VDD(VDD), .GND(GND), .A(G25), .Y(U376/a_13_43#));
	INVX1 X283 (.VDD(VDD), .GND(GND), .A(n223), .Y(n300));
	INVX1 X284 (.VDD(VDD), .GND(GND), .A(n295), .Y(n304));
	INVX1 X285 (.VDD(), .GND(), .A(n238), .Y());
	INVX1 X286 (.VDD(VDD), .GND(), .A(n234), .Y(n304));
	INVX1 X287 (.VDD(), .GND(), .A(n261), .Y());
	INVX1 X288 (.VDD(VDD), .GND(GND), .A(U379/a_13_43#), .Y(U379/a_18_54#));
	INVX1 X289 (.VDD(), .GND(), .A(n261), .Y());
	INVX1 X290 (.VDD(), .GND(), .A(U379/a_2_6#), .Y());
	INVX1 X291 (.VDD(), .GND(), .A(G24), .Y());
	INVX1 X292 (.VDD(VDD), .GND(GND), .A(G24), .Y(U379/a_13_43#));
	INVX1 X293 (.VDD(), .GND(), .A(n269), .Y());
	INVX1 X294 (.VDD(VDD), .GND(GND), .A(U380/a_13_43#), .Y(U380/a_18_54#));
	INVX1 X295 (.VDD(), .GND(), .A(n269), .Y());
	INVX1 X296 (.VDD(), .GND(), .A(U380/a_2_6#), .Y());
	INVX1 X297 (.VDD(), .GND(), .A(G23), .Y());
	INVX1 X298 (.VDD(VDD), .GND(GND), .A(G23), .Y(U380/a_13_43#));
	INVX1 X299 (.VDD(), .GND(), .A(n254), .Y());
	INVX1 X300 (.VDD(VDD), .GND(GND), .A(U381/a_13_43#), .Y(U381/a_18_54#));
	INVX1 X301 (.VDD(), .GND(), .A(n254), .Y());
	INVX1 X302 (.VDD(), .GND(), .A(U381/a_2_6#), .Y());
	INVX1 X303 (.VDD(), .GND(), .A(G22), .Y());
	INVX1 X304 (.VDD(VDD), .GND(GND), .A(G22), .Y(U381/a_13_43#));
	INVX1 X305 (.VDD(), .GND(), .A(n274), .Y());
	INVX1 X306 (.VDD(VDD), .GND(GND), .A(U382/a_13_43#), .Y(U382/a_18_54#));
	INVX1 X307 (.VDD(), .GND(), .A(n274), .Y());
	INVX1 X308 (.VDD(), .GND(), .A(U382/a_2_6#), .Y());
	INVX1 X309 (.VDD(), .GND(), .A(G21), .Y());
	INVX1 X310 (.VDD(VDD), .GND(GND), .A(G21), .Y(U382/a_13_43#));
	INVX1 X311 (.VDD(VDD), .GND(GND), .A(n224), .Y(n310));
	INVX1 X312 (.VDD(VDD), .GND(GND), .A(n294), .Y(n314));
	INVX1 X313 (.VDD(), .GND(), .A(n238), .Y());
	INVX1 X314 (.VDD(VDD), .GND(), .A(n235), .Y(n314));
	INVX1 X315 (.VDD(), .GND(), .A(n253), .Y());
	INVX1 X316 (.VDD(VDD), .GND(GND), .A(U385/a_13_43#), .Y(U385/a_18_54#));
	INVX1 X317 (.VDD(), .GND(), .A(n253), .Y());
	INVX1 X318 (.VDD(), .GND(), .A(U385/a_2_6#), .Y());
	INVX1 X319 (.VDD(), .GND(), .A(G20), .Y());
	INVX1 X320 (.VDD(VDD), .GND(GND), .A(G20), .Y(U385/a_13_43#));
	INVX1 X321 (.VDD(), .GND(), .A(n247), .Y());
	INVX1 X322 (.VDD(VDD), .GND(GND), .A(U386/a_13_43#), .Y(U386/a_18_54#));
	INVX1 X323 (.VDD(), .GND(), .A(n247), .Y());
	INVX1 X324 (.VDD(), .GND(), .A(U386/a_2_6#), .Y());
	INVX1 X325 (.VDD(), .GND(), .A(G19), .Y());
	INVX1 X326 (.VDD(VDD), .GND(GND), .A(G19), .Y(U386/a_13_43#));
	INVX1 X327 (.VDD(), .GND(), .A(n260), .Y());
	INVX1 X328 (.VDD(VDD), .GND(GND), .A(U387/a_13_43#), .Y(U387/a_18_54#));
	INVX1 X329 (.VDD(), .GND(), .A(n260), .Y());
	INVX1 X330 (.VDD(), .GND(), .A(U387/a_2_6#), .Y());
	INVX1 X331 (.VDD(), .GND(), .A(G18), .Y());
	INVX1 X332 (.VDD(VDD), .GND(GND), .A(G18), .Y(U387/a_13_43#));
	INVX1 X333 (.VDD(), .GND(), .A(n268), .Y());
	INVX1 X334 (.VDD(VDD), .GND(GND), .A(U388/a_13_43#), .Y(U388/a_18_54#));
	INVX1 X335 (.VDD(), .GND(), .A(n268), .Y());
	INVX1 X336 (.VDD(), .GND(), .A(U388/a_2_6#), .Y());
	INVX1 X337 (.VDD(), .GND(), .A(G17), .Y());
	INVX1 X338 (.VDD(VDD), .GND(GND), .A(G17), .Y(U388/a_13_43#));
	INVX1 X339 (.VDD(VDD), .GND(GND), .A(n225), .Y(n319));
	INVX1 X340 (.VDD(VDD), .GND(), .A(n297), .Y(n323));
	INVX1 X341 (.VDD(), .GND(), .A(n298), .Y());
	INVX1 X342 (.VDD(VDD), .GND(GND), .A(n324), .Y(n323));
	INVX1 X343 (.VDD(), .GND(GND), .A(n295), .Y(U427/a_9_6#));
	INVX1 X344 (.VDD(VDD), .GND(GND), .A(n295), .Y(U391/a_2_64#));
	INVX1 X345 (.VDD(), .GND(GND), .A(n294), .Y(n324));
	INVX1 X346 (.VDD(), .GND(GND), .A(n294), .Y(U430/a_9_6#));
	INVX1 X347 (.VDD(VDD), .GND(GND), .A(n327), .Y(n326));
	INVX1 X348 (.VDD(), .GND(), .A(n277), .Y());
	INVX1 X349 (.VDD(VDD), .GND(), .A(n329), .Y(n326));
	INVX1 X350 (.VDD(VDD), .GND(GND), .A(n330), .Y(n325));
	INVX1 X351 (.VDD(), .GND(), .A(n283), .Y());
	INVX1 X352 (.VDD(VDD), .GND(), .A(n332), .Y(n325));
	INVX1 X353 (.VDD(), .GND(), .A(n273), .Y());
	INVX1 X354 (.VDD(VDD), .GND(GND), .A(U394/a_13_43#), .Y(U394/a_18_54#));
	INVX1 X355 (.VDD(), .GND(), .A(n273), .Y());
	INVX1 X356 (.VDD(), .GND(), .A(U394/a_2_6#), .Y());
	INVX1 X357 (.VDD(), .GND(), .A(G16), .Y());
	INVX1 X358 (.VDD(VDD), .GND(GND), .A(G16), .Y(U394/a_13_43#));
	INVX1 X359 (.VDD(), .GND(), .A(n279), .Y());
	INVX1 X360 (.VDD(VDD), .GND(GND), .A(U395/a_13_43#), .Y(U395/a_18_54#));
	INVX1 X361 (.VDD(), .GND(), .A(n279), .Y());
	INVX1 X362 (.VDD(), .GND(), .A(U395/a_2_6#), .Y());
	INVX1 X363 (.VDD(), .GND(), .A(G15), .Y());
	INVX1 X364 (.VDD(VDD), .GND(GND), .A(G15), .Y(U395/a_13_43#));
	INVX1 X365 (.VDD(), .GND(), .A(n267), .Y());
	INVX1 X366 (.VDD(VDD), .GND(GND), .A(U396/a_13_43#), .Y(U396/a_18_54#));
	INVX1 X367 (.VDD(), .GND(), .A(n267), .Y());
	INVX1 X368 (.VDD(), .GND(), .A(U396/a_2_6#), .Y());
	INVX1 X369 (.VDD(), .GND(), .A(G14), .Y());
	INVX1 X370 (.VDD(VDD), .GND(GND), .A(G14), .Y(U396/a_13_43#));
	INVX1 X371 (.VDD(), .GND(), .A(n256), .Y());
	INVX1 X372 (.VDD(VDD), .GND(GND), .A(U397/a_12_41#), .Y(U397/a_18_54#));
	INVX1 X373 (.VDD(), .GND(), .A(U397/a_2_6#), .Y());
	INVX1 X374 (.VDD(), .GND(), .A(n256), .Y());
	INVX1 X375 (.VDD(), .GND(), .A(n339), .Y());
	INVX1 X376 (.VDD(VDD), .GND(GND), .A(n339), .Y(U397/a_12_41#));
	INVX1 X377 (.VDD(VDD), .GND(GND), .A(n226), .Y(n334));
	INVX1 X378 (.VDD(VDD), .GND(GND), .A(n327), .Y(n341));
	INVX1 X379 (.VDD(), .GND(), .A(n332), .Y());
	INVX1 X380 (.VDD(VDD), .GND(), .A(n342), .Y(n341));
	INVX1 X381 (.VDD(), .GND(GND), .A(n329), .Y(n342));
	INVX1 X382 (.VDD(VDD), .GND(), .A(n329), .Y(U400/a_2_64#));
	INVX1 X383 (.VDD(), .GND(), .A(n350), .Y());
	INVX1 X384 (.VDD(), .GND(), .A(n350), .Y());
	INVX1 X385 (.VDD(), .GND(GND), .A(n330), .Y(n342));
	INVX1 X386 (.VDD(), .GND(GND), .A(n330), .Y(U412/a_9_6#));
	INVX1 X387 (.VDD(), .GND(), .A(n266), .Y());
	INVX1 X388 (.VDD(VDD), .GND(GND), .A(U401/a_13_43#), .Y(U401/a_18_54#));
	INVX1 X389 (.VDD(), .GND(), .A(n266), .Y());
	INVX1 X390 (.VDD(), .GND(), .A(U401/a_2_6#), .Y());
	INVX1 X391 (.VDD(), .GND(), .A(G12), .Y());
	INVX1 X392 (.VDD(VDD), .GND(GND), .A(G12), .Y(U401/a_13_43#));
	INVX1 X393 (.VDD(), .GND(), .A(n259), .Y());
	INVX1 X394 (.VDD(VDD), .GND(GND), .A(U402/a_13_43#), .Y(U402/a_18_54#));
	INVX1 X395 (.VDD(), .GND(), .A(n259), .Y());
	INVX1 X396 (.VDD(), .GND(), .A(U402/a_2_6#), .Y());
	INVX1 X397 (.VDD(), .GND(), .A(G11), .Y());
	INVX1 X398 (.VDD(VDD), .GND(GND), .A(G11), .Y(U402/a_13_43#));
	INVX1 X399 (.VDD(), .GND(), .A(n241), .Y());
	INVX1 X400 (.VDD(VDD), .GND(GND), .A(U403/a_12_41#), .Y(U403/a_18_54#));
	INVX1 X401 (.VDD(), .GND(), .A(U403/a_2_6#), .Y());
	INVX1 X402 (.VDD(), .GND(), .A(n241), .Y());
	INVX1 X403 (.VDD(), .GND(), .A(n347), .Y());
	INVX1 X404 (.VDD(VDD), .GND(GND), .A(n347), .Y(U403/a_12_41#));
	INVX1 X405 (.VDD(), .GND(), .A(n252), .Y());
	INVX1 X406 (.VDD(VDD), .GND(GND), .A(U404/a_13_43#), .Y(U404/a_18_54#));
	INVX1 X407 (.VDD(), .GND(), .A(n252), .Y());
	INVX1 X408 (.VDD(), .GND(), .A(U404/a_2_6#), .Y());
	INVX1 X409 (.VDD(), .GND(), .A(G9), .Y());
	INVX1 X410 (.VDD(VDD), .GND(GND), .A(G9), .Y(U404/a_13_43#));
	INVX1 X411 (.VDD(VDD), .GND(GND), .A(n227), .Y(n344));
	INVX1 X412 (.VDD(VDD), .GND(GND), .A(n327), .Y(n349));
	INVX1 X413 (.VDD(), .GND(), .A(n239), .Y());
	INVX1 X414 (.VDD(VDD), .GND(), .A(n236), .Y(n349));
	INVX1 X415 (.VDD(), .GND(), .A(n258), .Y());
	INVX1 X416 (.VDD(VDD), .GND(GND), .A(U407/a_13_43#), .Y(U407/a_18_54#));
	INVX1 X417 (.VDD(), .GND(), .A(n258), .Y());
	INVX1 X418 (.VDD(), .GND(), .A(U407/a_2_6#), .Y());
	INVX1 X419 (.VDD(), .GND(), .A(G8), .Y());
	INVX1 X420 (.VDD(VDD), .GND(GND), .A(G8), .Y(U407/a_13_43#));
	INVX1 X421 (.VDD(), .GND(), .A(n265), .Y());
	INVX1 X422 (.VDD(VDD), .GND(GND), .A(U408/a_13_43#), .Y(U408/a_18_54#));
	INVX1 X423 (.VDD(), .GND(), .A(n265), .Y());
	INVX1 X424 (.VDD(), .GND(), .A(U408/a_2_6#), .Y());
	INVX1 X425 (.VDD(), .GND(), .A(G7), .Y());
	INVX1 X426 (.VDD(VDD), .GND(GND), .A(G7), .Y(U408/a_13_43#));
	INVX1 X427 (.VDD(), .GND(), .A(n251), .Y());
	INVX1 X428 (.VDD(VDD), .GND(GND), .A(U409/a_13_43#), .Y(U409/a_18_54#));
	INVX1 X429 (.VDD(), .GND(), .A(n251), .Y());
	INVX1 X430 (.VDD(), .GND(), .A(U409/a_2_6#), .Y());
	INVX1 X431 (.VDD(), .GND(), .A(G6), .Y());
	INVX1 X432 (.VDD(VDD), .GND(GND), .A(G6), .Y(U409/a_13_43#));
	INVX1 X433 (.VDD(), .GND(), .A(n240), .Y());
	INVX1 X434 (.VDD(VDD), .GND(GND), .A(U410/a_12_41#), .Y(U410/a_18_54#));
	INVX1 X435 (.VDD(), .GND(), .A(U410/a_2_6#), .Y());
	INVX1 X436 (.VDD(), .GND(), .A(n240), .Y());
	INVX1 X437 (.VDD(), .GND(), .A(n357), .Y());
	INVX1 X438 (.VDD(VDD), .GND(GND), .A(n357), .Y(U410/a_12_41#));
	INVX1 X439 (.VDD(VDD), .GND(GND), .A(n228), .Y(n353));
	INVX1 X440 (.VDD(VDD), .GND(), .A(n330), .Y(n358));
	INVX1 X441 (.VDD(), .GND(), .A(n239), .Y());
	INVX1 X442 (.VDD(), .GND(), .A(n250), .Y());
	INVX1 X443 (.VDD(VDD), .GND(GND), .A(U413/a_13_43#), .Y(U413/a_18_54#));
	INVX1 X444 (.VDD(), .GND(), .A(n250), .Y());
	INVX1 X445 (.VDD(), .GND(), .A(U413/a_2_6#), .Y());
	INVX1 X446 (.VDD(), .GND(), .A(G4), .Y());
	INVX1 X447 (.VDD(VDD), .GND(GND), .A(G4), .Y(U413/a_13_43#));
	INVX1 X448 (.VDD(), .GND(), .A(n246), .Y());
	INVX1 X449 (.VDD(VDD), .GND(GND), .A(U414/a_13_43#), .Y(U414/a_18_54#));
	INVX1 X450 (.VDD(), .GND(), .A(n246), .Y());
	INVX1 X451 (.VDD(), .GND(), .A(U414/a_2_6#), .Y());
	INVX1 X452 (.VDD(), .GND(), .A(G3), .Y());
	INVX1 X453 (.VDD(VDD), .GND(GND), .A(G3), .Y(U414/a_13_43#));
	INVX1 X454 (.VDD(), .GND(), .A(n278), .Y());
	INVX1 X455 (.VDD(VDD), .GND(GND), .A(U415/a_13_43#), .Y(U415/a_18_54#));
	INVX1 X456 (.VDD(), .GND(), .A(n278), .Y());
	INVX1 X457 (.VDD(), .GND(), .A(U415/a_2_6#), .Y());
	INVX1 X458 (.VDD(), .GND(), .A(G2), .Y());
	INVX1 X459 (.VDD(VDD), .GND(GND), .A(G2), .Y(U415/a_13_43#));
	INVX1 X460 (.VDD(), .GND(), .A(n272), .Y());
	INVX1 X461 (.VDD(VDD), .GND(GND), .A(U416/a_13_43#), .Y(U416/a_18_54#));
	INVX1 X462 (.VDD(), .GND(), .A(n272), .Y());
	INVX1 X463 (.VDD(), .GND(), .A(U416/a_2_6#), .Y());
	INVX1 X464 (.VDD(), .GND(), .A(G1), .Y());
	INVX1 X465 (.VDD(VDD), .GND(GND), .A(G1), .Y(U416/a_13_43#));
	INVX1 X466 (.VDD(VDD), .GND(GND), .A(n229), .Y(n361));
	INVX1 X467 (.VDD(VDD), .GND(GND), .A(n330), .Y(n365));
	INVX1 X468 (.VDD(), .GND(), .A(n329), .Y());
	INVX1 X469 (.VDD(VDD), .GND(GND), .A(n366), .Y(n365));
	INVX1 X470 (.VDD(), .GND(GND), .A(n327), .Y(n327));
	INVX1 X471 (.VDD(), .GND(GND), .A(n332), .Y(n366));
	INVX1 X472 (.VDD(), .GND(GND), .A(n332), .Y(n332));
	INVX1 X473 (.VDD(VDD), .GND(), .A(n288), .Y(n332));
	INVX1 X474 (.VDD(), .GND(), .A(n367), .Y());
	INVX1 X475 (.VDD(VDD), .GND(GND), .A(U421/a_12_41#), .Y(U421/a_18_54#));
	INVX1 X476 (.VDD(), .GND(), .A(U421/a_2_6#), .Y());
	INVX1 X477 (.VDD(), .GND(), .A(n367), .Y());
	INVX1 X478 (.VDD(), .GND(), .A(n368), .Y());
	INVX1 X479 (.VDD(VDD), .GND(GND), .A(n368), .Y(U421/a_12_41#));
	INVX1 X480 (.VDD(), .GND(), .A(n369), .Y());
	INVX1 X481 (.VDD(VDD), .GND(GND), .A(U422/a_13_43#), .Y(U422/a_18_54#));
	INVX1 X482 (.VDD(), .GND(), .A(n369), .Y());
	INVX1 X483 (.VDD(), .GND(), .A(U422/a_2_6#), .Y());
	INVX1 X484 (.VDD(), .GND(), .A(n370), .Y());
	INVX1 X485 (.VDD(VDD), .GND(GND), .A(n370), .Y(U422/a_13_43#));
	INVX1 X486 (.VDD(), .GND(), .A(G23), .Y());
	INVX1 X487 (.VDD(VDD), .GND(GND), .A(U423/a_13_43#), .Y(U423/a_18_54#));
	INVX1 X488 (.VDD(), .GND(), .A(G23), .Y());
	INVX1 X489 (.VDD(), .GND(), .A(U423/a_2_6#), .Y());
	INVX1 X490 (.VDD(), .GND(), .A(G19), .Y());
	INVX1 X491 (.VDD(VDD), .GND(GND), .A(G19), .Y(U423/a_13_43#));
	INVX1 X492 (.VDD(), .GND(), .A(G31), .Y());
	INVX1 X493 (.VDD(VDD), .GND(GND), .A(U424/a_13_43#), .Y(U424/a_18_54#));
	INVX1 X494 (.VDD(), .GND(), .A(G31), .Y());
	INVX1 X495 (.VDD(), .GND(), .A(U424/a_2_6#), .Y());
	INVX1 X496 (.VDD(), .GND(), .A(G27), .Y());
	INVX1 X497 (.VDD(VDD), .GND(GND), .A(G27), .Y(U424/a_13_43#));
	INVX1 X498 (.VDD(), .GND(), .A(n371), .Y());
	INVX1 X499 (.VDD(VDD), .GND(GND), .A(U425/a_13_43#), .Y(U425/a_18_54#));
	INVX1 X500 (.VDD(), .GND(), .A(n371), .Y());
	INVX1 X501 (.VDD(), .GND(), .A(n372), .Y());
	INVX1 X502 (.VDD(VDD), .GND(GND), .A(n372), .Y(U425/a_13_43#));
	INVX1 X503 (.VDD(), .GND(), .A(n248), .Y());
	INVX1 X504 (.VDD(VDD), .GND(GND), .A(U426/a_13_43#), .Y(U426/a_18_54#));
	INVX1 X505 (.VDD(), .GND(), .A(n248), .Y());
	INVX1 X506 (.VDD(), .GND(), .A(U426/a_2_6#), .Y());
	INVX1 X507 (.VDD(), .GND(), .A(n374), .Y());
	INVX1 X508 (.VDD(VDD), .GND(GND), .A(n374), .Y(U426/a_13_43#));
	INVX1 X509 (.VDD(), .GND(), .A(n276), .Y());
	INVX1 X510 (.VDD(VDD), .GND(GND), .A(n298), .Y(n376));
	INVX1 X511 (.VDD(VDD), .GND(), .A(n307), .Y(n298));
	INVX1 X512 (.VDD(VDD), .GND(), .A(n340), .Y(n295));
	INVX1 X513 (.VDD(VDD), .GND(), .A(n294), .Y(n375));
	INVX1 X514 (.VDD(), .GND(), .A(n282), .Y());
	INVX1 X515 (.VDD(VDD), .GND(GND), .A(n297), .Y(n375));
	INVX1 X516 (.VDD(VDD), .GND(), .A(n316), .Y(n297));
	INVX1 X517 (.VDD(), .GND(), .A(n377), .Y());
	INVX1 X518 (.VDD(VDD), .GND(GND), .A(U432/a_12_41#), .Y(U432/a_18_54#));
	INVX1 X519 (.VDD(), .GND(), .A(U432/a_2_6#), .Y());
	INVX1 X520 (.VDD(), .GND(), .A(n377), .Y());
	INVX1 X521 (.VDD(), .GND(), .A(n378), .Y());
	INVX1 X522 (.VDD(VDD), .GND(GND), .A(n378), .Y(U432/a_12_41#));
	INVX1 X523 (.VDD(), .GND(), .A(n379), .Y());
	INVX1 X524 (.VDD(VDD), .GND(GND), .A(U433/a_13_43#), .Y(U433/a_18_54#));
	INVX1 X525 (.VDD(), .GND(), .A(n379), .Y());
	INVX1 X526 (.VDD(), .GND(), .A(U433/a_2_6#), .Y());
	INVX1 X527 (.VDD(), .GND(), .A(n380), .Y());
	INVX1 X528 (.VDD(VDD), .GND(GND), .A(n380), .Y(U433/a_13_43#));
	INVX1 X529 (.VDD(), .GND(), .A(G14), .Y());
	INVX1 X530 (.VDD(VDD), .GND(GND), .A(U434/a_12_41#), .Y(U434/a_18_54#));
	INVX1 X531 (.VDD(), .GND(), .A(U434/a_2_6#), .Y());
	INVX1 X532 (.VDD(), .GND(), .A(G14), .Y());
	INVX1 X533 (.VDD(), .GND(), .A(n347), .Y());
	INVX1 X534 (.VDD(VDD), .GND(GND), .A(n347), .Y(U434/a_12_41#));
	INVX1 X535 (.VDD(VDD), .GND(GND), .A(G10), .Y(n347));
	INVX1 X536 (.VDD(), .GND(), .A(G6), .Y());
	INVX1 X537 (.VDD(VDD), .GND(GND), .A(U436/a_13_43#), .Y(U436/a_18_54#));
	INVX1 X538 (.VDD(), .GND(), .A(G6), .Y());
	INVX1 X539 (.VDD(), .GND(), .A(U436/a_2_6#), .Y());
	INVX1 X540 (.VDD(), .GND(), .A(G2), .Y());
	INVX1 X541 (.VDD(VDD), .GND(GND), .A(G2), .Y(U436/a_13_43#));
	INVX1 X542 (.VDD(), .GND(), .A(n381), .Y());
	INVX1 X543 (.VDD(VDD), .GND(GND), .A(U437/a_13_43#), .Y(U437/a_18_54#));
	INVX1 X544 (.VDD(), .GND(), .A(n381), .Y());
	INVX1 X545 (.VDD(), .GND(), .A(n382), .Y());
	INVX1 X546 (.VDD(VDD), .GND(GND), .A(n382), .Y(U437/a_13_43#));
	INVX1 X547 (.VDD(), .GND(), .A(n257), .Y());
	INVX1 X548 (.VDD(VDD), .GND(GND), .A(U438/a_13_43#), .Y(U438/a_18_54#));
	INVX1 X549 (.VDD(), .GND(), .A(n257), .Y());
	INVX1 X550 (.VDD(), .GND(), .A(U438/a_2_6#), .Y());
	INVX1 X551 (.VDD(), .GND(), .A(n384), .Y());
	INVX1 X552 (.VDD(VDD), .GND(GND), .A(n384), .Y(U438/a_13_43#));
	INVX1 X553 (.VDD(), .GND(), .A(n385), .Y());
	INVX1 X554 (.VDD(VDD), .GND(GND), .A(U439/a_12_41#), .Y(U439/a_18_54#));
	INVX1 X555 (.VDD(), .GND(), .A(U439/a_2_6#), .Y());
	INVX1 X556 (.VDD(), .GND(), .A(n385), .Y());
	INVX1 X557 (.VDD(), .GND(), .A(n386), .Y());
	INVX1 X558 (.VDD(VDD), .GND(GND), .A(n386), .Y(U439/a_12_41#));
	INVX1 X559 (.VDD(), .GND(), .A(n387), .Y());
	INVX1 X560 (.VDD(VDD), .GND(GND), .A(U440/a_13_43#), .Y(U440/a_18_54#));
	INVX1 X561 (.VDD(), .GND(), .A(n387), .Y());
	INVX1 X562 (.VDD(), .GND(), .A(U440/a_2_6#), .Y());
	INVX1 X563 (.VDD(), .GND(), .A(n388), .Y());
	INVX1 X564 (.VDD(VDD), .GND(GND), .A(n388), .Y(U440/a_13_43#));
	INVX1 X565 (.VDD(), .GND(), .A(G16), .Y());
	INVX1 X566 (.VDD(VDD), .GND(GND), .A(U441/a_13_43#), .Y(U441/a_18_54#));
	INVX1 X567 (.VDD(), .GND(), .A(G16), .Y());
	INVX1 X568 (.VDD(), .GND(), .A(U441/a_2_6#), .Y());
	INVX1 X569 (.VDD(), .GND(), .A(G12), .Y());
	INVX1 X570 (.VDD(VDD), .GND(GND), .A(G12), .Y(U441/a_13_43#));
	INVX1 X571 (.VDD(), .GND(), .A(G8), .Y());
	INVX1 X572 (.VDD(VDD), .GND(GND), .A(U442/a_13_43#), .Y(U442/a_18_54#));
	INVX1 X573 (.VDD(), .GND(), .A(G8), .Y());
	INVX1 X574 (.VDD(), .GND(), .A(U442/a_2_6#), .Y());
	INVX1 X575 (.VDD(), .GND(), .A(G4), .Y());
	INVX1 X576 (.VDD(VDD), .GND(GND), .A(G4), .Y(U442/a_13_43#));
	INVX1 X577 (.VDD(), .GND(), .A(n389), .Y());
	INVX1 X578 (.VDD(VDD), .GND(GND), .A(U443/a_13_43#), .Y(U443/a_18_54#));
	INVX1 X579 (.VDD(), .GND(), .A(n389), .Y());
	INVX1 X580 (.VDD(), .GND(), .A(n390), .Y());
	INVX1 X581 (.VDD(VDD), .GND(GND), .A(n390), .Y(U443/a_13_43#));
	INVX1 X582 (.VDD(), .GND(), .A(n242), .Y());
	INVX1 X583 (.VDD(VDD), .GND(GND), .A(U444/a_13_43#), .Y(U444/a_18_54#));
	INVX1 X584 (.VDD(), .GND(), .A(n242), .Y());
	INVX1 X585 (.VDD(), .GND(), .A(U444/a_2_6#), .Y());
	INVX1 X586 (.VDD(), .GND(), .A(n384), .Y());
	INVX1 X587 (.VDD(VDD), .GND(GND), .A(n384), .Y(U444/a_13_43#));
	INVX1 X588 (.VDD(), .GND(), .A(n392), .Y());
	INVX1 X589 (.VDD(VDD), .GND(GND), .A(U445/a_12_41#), .Y(U445/a_18_54#));
	INVX1 X590 (.VDD(), .GND(), .A(U445/a_2_6#), .Y());
	INVX1 X591 (.VDD(), .GND(), .A(n392), .Y());
	INVX1 X592 (.VDD(), .GND(), .A(n393), .Y());
	INVX1 X593 (.VDD(VDD), .GND(GND), .A(n393), .Y(U445/a_12_41#));
	INVX1 X594 (.VDD(), .GND(), .A(G32), .Y());
	INVX1 X595 (.VDD(VDD), .GND(GND), .A(U446/a_13_43#), .Y(U446/a_18_54#));
	INVX1 X596 (.VDD(), .GND(), .A(G32), .Y());
	INVX1 X597 (.VDD(), .GND(), .A(U446/a_2_6#), .Y());
	INVX1 X598 (.VDD(), .GND(), .A(G31), .Y());
	INVX1 X599 (.VDD(VDD), .GND(GND), .A(G31), .Y(U446/a_13_43#));
	INVX1 X600 (.VDD(), .GND(), .A(G29), .Y());
	INVX1 X601 (.VDD(VDD), .GND(GND), .A(U447/a_12_41#), .Y(U447/a_18_54#));
	INVX1 X602 (.VDD(), .GND(), .A(U447/a_2_6#), .Y());
	INVX1 X603 (.VDD(), .GND(), .A(G29), .Y());
	INVX1 X604 (.VDD(), .GND(), .A(G30), .Y());
	INVX1 X605 (.VDD(VDD), .GND(GND), .A(G30), .Y(U447/a_12_41#));
	INVX1 X606 (.VDD(), .GND(), .A(n394), .Y());
	INVX1 X607 (.VDD(VDD), .GND(GND), .A(U448/a_12_41#), .Y(U448/a_18_54#));
	INVX1 X608 (.VDD(), .GND(), .A(U448/a_2_6#), .Y());
	INVX1 X609 (.VDD(), .GND(), .A(n394), .Y());
	INVX1 X610 (.VDD(), .GND(), .A(n395), .Y());
	INVX1 X611 (.VDD(VDD), .GND(GND), .A(n395), .Y(U448/a_12_41#));
	INVX1 X612 (.VDD(), .GND(), .A(n396), .Y());
	INVX1 X613 (.VDD(VDD), .GND(GND), .A(U449/a_13_43#), .Y(U449/a_18_54#));
	INVX1 X614 (.VDD(), .GND(), .A(n396), .Y());
	INVX1 X615 (.VDD(), .GND(), .A(U449/a_2_6#), .Y());
	INVX1 X616 (.VDD(), .GND(), .A(n397), .Y());
	INVX1 X617 (.VDD(VDD), .GND(GND), .A(n397), .Y(U449/a_13_43#));
	INVX1 X618 (.VDD(), .GND(), .A(n339), .Y());
	INVX1 X619 (.VDD(VDD), .GND(GND), .A(U450/a_12_41#), .Y(U450/a_18_54#));
	INVX1 X620 (.VDD(), .GND(), .A(U450/a_2_6#), .Y());
	INVX1 X621 (.VDD(), .GND(), .A(n339), .Y());
	INVX1 X622 (.VDD(), .GND(), .A(G1), .Y());
	INVX1 X623 (.VDD(VDD), .GND(GND), .A(G1), .Y(U450/a_12_41#));
	INVX1 X624 (.VDD(VDD), .GND(GND), .A(G13), .Y(n339));
	INVX1 X625 (.VDD(), .GND(), .A(G9), .Y());
	INVX1 X626 (.VDD(VDD), .GND(GND), .A(U452/a_12_41#), .Y(U452/a_18_54#));
	INVX1 X627 (.VDD(), .GND(), .A(U452/a_2_6#), .Y());
	INVX1 X628 (.VDD(), .GND(), .A(G9), .Y());
	INVX1 X629 (.VDD(), .GND(), .A(n357), .Y());
	INVX1 X630 (.VDD(VDD), .GND(GND), .A(n357), .Y(U452/a_12_41#));
	INVX1 X631 (.VDD(VDD), .GND(GND), .A(G5), .Y(n357));
	INVX1 X632 (.VDD(), .GND(), .A(n398), .Y());
	INVX1 X633 (.VDD(VDD), .GND(GND), .A(U454/a_13_43#), .Y(U454/a_18_54#));
	INVX1 X634 (.VDD(), .GND(), .A(n398), .Y());
	INVX1 X635 (.VDD(), .GND(), .A(n399), .Y());
	INVX1 X636 (.VDD(VDD), .GND(GND), .A(n399), .Y(U454/a_13_43#));
	INVX1 X637 (.VDD(), .GND(), .A(n264), .Y());
	INVX1 X638 (.VDD(VDD), .GND(GND), .A(U455/a_13_43#), .Y(U455/a_18_54#));
	INVX1 X639 (.VDD(), .GND(), .A(n264), .Y());
	INVX1 X640 (.VDD(), .GND(), .A(U455/a_2_6#), .Y());
	INVX1 X641 (.VDD(), .GND(), .A(n390), .Y());
	INVX1 X642 (.VDD(VDD), .GND(GND), .A(n390), .Y(U455/a_13_43#));
	INVX1 X643 (.VDD(), .GND(), .A(n401), .Y());
	INVX1 X644 (.VDD(VDD), .GND(GND), .A(U456/a_12_41#), .Y(U456/a_18_54#));
	INVX1 X645 (.VDD(), .GND(), .A(U456/a_2_6#), .Y());
	INVX1 X646 (.VDD(), .GND(), .A(n401), .Y());
	INVX1 X647 (.VDD(), .GND(), .A(n402), .Y());
	INVX1 X648 (.VDD(VDD), .GND(GND), .A(n402), .Y(U456/a_12_41#));
	INVX1 X649 (.VDD(), .GND(), .A(G24), .Y());
	INVX1 X650 (.VDD(VDD), .GND(GND), .A(U457/a_13_43#), .Y(U457/a_18_54#));
	INVX1 X651 (.VDD(), .GND(), .A(G24), .Y());
	INVX1 X652 (.VDD(), .GND(), .A(U457/a_2_6#), .Y());
	INVX1 X653 (.VDD(), .GND(), .A(G23), .Y());
	INVX1 X654 (.VDD(VDD), .GND(GND), .A(G23), .Y(U457/a_13_43#));
	INVX1 X655 (.VDD(), .GND(), .A(G21), .Y());
	INVX1 X656 (.VDD(VDD), .GND(GND), .A(U458/a_12_41#), .Y(U458/a_18_54#));
	INVX1 X657 (.VDD(), .GND(), .A(U458/a_2_6#), .Y());
	INVX1 X658 (.VDD(), .GND(), .A(G21), .Y());
	INVX1 X659 (.VDD(), .GND(), .A(G22), .Y());
	INVX1 X660 (.VDD(VDD), .GND(GND), .A(G22), .Y(U458/a_12_41#));
	INVX1 X661 (.VDD(VDD), .GND(GND), .A(n336), .Y(n294));
	INVX1 X662 (.VDD(), .GND(), .A(n403), .Y());
	INVX1 X663 (.VDD(VDD), .GND(GND), .A(U460/a_12_41#), .Y(U460/a_18_54#));
	INVX1 X664 (.VDD(), .GND(), .A(U460/a_2_6#), .Y());
	INVX1 X665 (.VDD(), .GND(), .A(n403), .Y());
	INVX1 X666 (.VDD(), .GND(), .A(n404), .Y());
	INVX1 X667 (.VDD(VDD), .GND(GND), .A(n404), .Y(U460/a_12_41#));
	INVX1 X668 (.VDD(), .GND(), .A(n405), .Y());
	INVX1 X669 (.VDD(VDD), .GND(GND), .A(U461/a_13_43#), .Y(U461/a_18_54#));
	INVX1 X670 (.VDD(), .GND(), .A(n405), .Y());
	INVX1 X671 (.VDD(), .GND(), .A(U461/a_2_6#), .Y());
	INVX1 X672 (.VDD(), .GND(), .A(n406), .Y());
	INVX1 X673 (.VDD(VDD), .GND(GND), .A(n406), .Y(U461/a_13_43#));
	INVX1 X674 (.VDD(), .GND(), .A(G15), .Y());
	INVX1 X675 (.VDD(VDD), .GND(GND), .A(U462/a_13_43#), .Y(U462/a_18_54#));
	INVX1 X676 (.VDD(), .GND(), .A(G15), .Y());
	INVX1 X677 (.VDD(), .GND(), .A(U462/a_2_6#), .Y());
	INVX1 X678 (.VDD(), .GND(), .A(G11), .Y());
	INVX1 X679 (.VDD(VDD), .GND(GND), .A(G11), .Y(U462/a_13_43#));
	INVX1 X680 (.VDD(), .GND(), .A(G7), .Y());
	INVX1 X681 (.VDD(VDD), .GND(GND), .A(U463/a_13_43#), .Y(U463/a_18_54#));
	INVX1 X682 (.VDD(), .GND(), .A(G7), .Y());
	INVX1 X683 (.VDD(), .GND(), .A(U463/a_2_6#), .Y());
	INVX1 X684 (.VDD(), .GND(), .A(G3), .Y());
	INVX1 X685 (.VDD(VDD), .GND(GND), .A(G3), .Y(U463/a_13_43#));
	INVX1 X686 (.VDD(), .GND(), .A(n407), .Y());
	INVX1 X687 (.VDD(VDD), .GND(GND), .A(U464/a_13_43#), .Y(U464/a_18_54#));
	INVX1 X688 (.VDD(), .GND(), .A(n407), .Y());
	INVX1 X689 (.VDD(), .GND(), .A(U464/a_2_6#), .Y());
	INVX1 X690 (.VDD(), .GND(), .A(n399), .Y());
	INVX1 X691 (.VDD(VDD), .GND(GND), .A(n399), .Y(U464/a_13_43#));
	INVX1 X692 (.VDD(), .GND(), .A(n408), .Y());
	INVX1 X693 (.VDD(VDD), .GND(GND), .A(U465/a_12_41#), .Y(U465/a_18_54#));
	INVX1 X694 (.VDD(), .GND(), .A(U465/a_2_6#), .Y());
	INVX1 X695 (.VDD(), .GND(), .A(n408), .Y());
	INVX1 X696 (.VDD(), .GND(), .A(n409), .Y());
	INVX1 X697 (.VDD(VDD), .GND(GND), .A(n409), .Y(U465/a_12_41#));
	INVX1 X698 (.VDD(), .GND(), .A(G20), .Y());
	INVX1 X699 (.VDD(VDD), .GND(GND), .A(U466/a_13_43#), .Y(U466/a_18_54#));
	INVX1 X700 (.VDD(), .GND(), .A(G20), .Y());
	INVX1 X701 (.VDD(), .GND(), .A(U466/a_2_6#), .Y());
	INVX1 X702 (.VDD(), .GND(), .A(G19), .Y());
	INVX1 X703 (.VDD(VDD), .GND(GND), .A(G19), .Y(U466/a_13_43#));
	INVX1 X704 (.VDD(), .GND(), .A(G17), .Y());
	INVX1 X705 (.VDD(VDD), .GND(GND), .A(U467/a_12_41#), .Y(U467/a_18_54#));
	INVX1 X706 (.VDD(), .GND(), .A(U467/a_2_6#), .Y());
	INVX1 X707 (.VDD(), .GND(), .A(G17), .Y());
	INVX1 X708 (.VDD(), .GND(), .A(G18), .Y());
	INVX1 X709 (.VDD(VDD), .GND(GND), .A(G18), .Y(U467/a_12_41#));
	INVX1 X710 (.VDD(), .GND(), .A(n249), .Y());
	INVX1 X711 (.VDD(VDD), .GND(GND), .A(U468/a_13_43#), .Y(U468/a_18_54#));
	INVX1 X712 (.VDD(), .GND(), .A(n249), .Y());
	INVX1 X713 (.VDD(), .GND(), .A(U468/a_2_6#), .Y());
	INVX1 X714 (.VDD(), .GND(), .A(n382), .Y());
	INVX1 X715 (.VDD(VDD), .GND(GND), .A(n382), .Y(U468/a_13_43#));
	INVX1 X716 (.VDD(), .GND(), .A(n411), .Y());
	INVX1 X717 (.VDD(VDD), .GND(GND), .A(U469/a_12_41#), .Y(U469/a_18_54#));
	INVX1 X718 (.VDD(), .GND(), .A(U469/a_2_6#), .Y());
	INVX1 X719 (.VDD(), .GND(), .A(n411), .Y());
	INVX1 X720 (.VDD(), .GND(), .A(n412), .Y());
	INVX1 X721 (.VDD(VDD), .GND(GND), .A(n412), .Y(U469/a_12_41#));
	INVX1 X722 (.VDD(), .GND(), .A(G28), .Y());
	INVX1 X723 (.VDD(VDD), .GND(GND), .A(U470/a_13_43#), .Y(U470/a_18_54#));
	INVX1 X724 (.VDD(), .GND(), .A(G28), .Y());
	INVX1 X725 (.VDD(), .GND(), .A(U470/a_2_6#), .Y());
	INVX1 X726 (.VDD(), .GND(), .A(G27), .Y());
	INVX1 X727 (.VDD(VDD), .GND(GND), .A(G27), .Y(U470/a_13_43#));
	INVX1 X728 (.VDD(), .GND(), .A(G25), .Y());
	INVX1 X729 (.VDD(VDD), .GND(GND), .A(U471/a_12_41#), .Y(U471/a_18_54#));
	INVX1 X730 (.VDD(), .GND(), .A(U471/a_2_6#), .Y());
	INVX1 X731 (.VDD(), .GND(), .A(G25), .Y());
	INVX1 X732 (.VDD(), .GND(), .A(G26), .Y());
	INVX1 X733 (.VDD(VDD), .GND(GND), .A(G26), .Y(U471/a_12_41#));
	INVX1 X734 (.VDD(VDD), .GND(), .A(n292), .Y(n327));
	INVX1 X735 (.VDD(), .GND(), .A(n413), .Y());
	INVX1 X736 (.VDD(VDD), .GND(GND), .A(U473/a_12_41#), .Y(U473/a_18_54#));
	INVX1 X737 (.VDD(), .GND(), .A(U473/a_2_6#), .Y());
	INVX1 X738 (.VDD(), .GND(), .A(n413), .Y());
	INVX1 X739 (.VDD(), .GND(), .A(n414), .Y());
	INVX1 X740 (.VDD(VDD), .GND(GND), .A(n414), .Y(U473/a_12_41#));
	INVX1 X741 (.VDD(), .GND(), .A(n415), .Y());
	INVX1 X742 (.VDD(VDD), .GND(GND), .A(U474/a_13_43#), .Y(U474/a_18_54#));
	INVX1 X743 (.VDD(), .GND(), .A(n415), .Y());
	INVX1 X744 (.VDD(), .GND(), .A(U474/a_2_6#), .Y());
	INVX1 X745 (.VDD(), .GND(), .A(n416), .Y());
	INVX1 X746 (.VDD(VDD), .GND(GND), .A(n416), .Y(U474/a_13_43#));
	INVX1 X747 (.VDD(), .GND(), .A(G21), .Y());
	INVX1 X748 (.VDD(VDD), .GND(GND), .A(U475/a_13_43#), .Y(U475/a_18_54#));
	INVX1 X749 (.VDD(), .GND(), .A(G21), .Y());
	INVX1 X750 (.VDD(), .GND(), .A(U475/a_2_6#), .Y());
	INVX1 X751 (.VDD(), .GND(), .A(G17), .Y());
	INVX1 X752 (.VDD(VDD), .GND(GND), .A(G17), .Y(U475/a_13_43#));
	INVX1 X753 (.VDD(), .GND(), .A(G29), .Y());
	INVX1 X754 (.VDD(VDD), .GND(GND), .A(U476/a_13_43#), .Y(U476/a_18_54#));
	INVX1 X755 (.VDD(), .GND(), .A(G29), .Y());
	INVX1 X756 (.VDD(), .GND(), .A(U476/a_2_6#), .Y());
	INVX1 X757 (.VDD(), .GND(), .A(G25), .Y());
	INVX1 X758 (.VDD(VDD), .GND(GND), .A(G25), .Y(U476/a_13_43#));
	INVX1 X759 (.VDD(), .GND(), .A(n417), .Y());
	INVX1 X760 (.VDD(VDD), .GND(GND), .A(U477/a_13_43#), .Y(U477/a_18_54#));
	INVX1 X761 (.VDD(), .GND(), .A(n417), .Y());
	INVX1 X762 (.VDD(), .GND(), .A(n372), .Y());
	INVX1 X763 (.VDD(VDD), .GND(GND), .A(n372), .Y(U477/a_13_43#));
	INVX1 X764 (.VDD(), .GND(), .A(n418), .Y());
	INVX1 X765 (.VDD(VDD), .GND(GND), .A(U478/a_12_41#), .Y(U478/a_18_54#));
	INVX1 X766 (.VDD(), .GND(), .A(U478/a_2_6#), .Y());
	INVX1 X767 (.VDD(), .GND(), .A(n418), .Y());
	INVX1 X768 (.VDD(), .GND(), .A(n419), .Y());
	INVX1 X769 (.VDD(VDD), .GND(GND), .A(n419), .Y(U478/a_12_41#));
	INVX1 X770 (.VDD(), .GND(), .A(G4), .Y());
	INVX1 X771 (.VDD(VDD), .GND(GND), .A(U479/a_13_43#), .Y(U479/a_18_54#));
	INVX1 X772 (.VDD(), .GND(), .A(G4), .Y());
	INVX1 X773 (.VDD(), .GND(), .A(U479/a_2_6#), .Y());
	INVX1 X774 (.VDD(), .GND(), .A(G3), .Y());
	INVX1 X775 (.VDD(VDD), .GND(GND), .A(G3), .Y(U479/a_13_43#));
	INVX1 X776 (.VDD(), .GND(), .A(G1), .Y());
	INVX1 X777 (.VDD(VDD), .GND(GND), .A(U480/a_12_41#), .Y(U480/a_18_54#));
	INVX1 X778 (.VDD(), .GND(), .A(U480/a_2_6#), .Y());
	INVX1 X779 (.VDD(), .GND(), .A(G1), .Y());
	INVX1 X780 (.VDD(), .GND(), .A(G2), .Y());
	INVX1 X781 (.VDD(VDD), .GND(GND), .A(G2), .Y(U480/a_12_41#));
	INVX1 X782 (.VDD(), .GND(), .A(n244), .Y());
	INVX1 X783 (.VDD(VDD), .GND(GND), .A(U481/a_13_43#), .Y(U481/a_18_54#));
	INVX1 X784 (.VDD(), .GND(), .A(n244), .Y());
	INVX1 X785 (.VDD(), .GND(), .A(U481/a_2_6#), .Y());
	INVX1 X786 (.VDD(), .GND(), .A(n421), .Y());
	INVX1 X787 (.VDD(VDD), .GND(GND), .A(n421), .Y(U481/a_13_43#));
	INVX1 X788 (.VDD(VDD), .GND(GND), .A(n286), .Y(n329));
	INVX1 X789 (.VDD(), .GND(), .A(n422), .Y());
	INVX1 X790 (.VDD(VDD), .GND(GND), .A(U483/a_12_41#), .Y(U483/a_18_54#));
	INVX1 X791 (.VDD(), .GND(), .A(U483/a_2_6#), .Y());
	INVX1 X792 (.VDD(), .GND(), .A(n422), .Y());
	INVX1 X793 (.VDD(), .GND(), .A(n423), .Y());
	INVX1 X794 (.VDD(VDD), .GND(GND), .A(n423), .Y(U483/a_12_41#));
	INVX1 X795 (.VDD(), .GND(), .A(n424), .Y());
	INVX1 X796 (.VDD(VDD), .GND(GND), .A(U484/a_13_43#), .Y(U484/a_18_54#));
	INVX1 X797 (.VDD(), .GND(), .A(n424), .Y());
	INVX1 X798 (.VDD(), .GND(), .A(U484/a_2_6#), .Y());
	INVX1 X799 (.VDD(), .GND(), .A(n425), .Y());
	INVX1 X800 (.VDD(VDD), .GND(GND), .A(n425), .Y(U484/a_13_43#));
	INVX1 X801 (.VDD(), .GND(), .A(G24), .Y());
	INVX1 X802 (.VDD(VDD), .GND(GND), .A(U485/a_13_43#), .Y(U485/a_18_54#));
	INVX1 X803 (.VDD(), .GND(), .A(G24), .Y());
	INVX1 X804 (.VDD(), .GND(), .A(U485/a_2_6#), .Y());
	INVX1 X805 (.VDD(), .GND(), .A(G20), .Y());
	INVX1 X806 (.VDD(VDD), .GND(GND), .A(G20), .Y(U485/a_13_43#));
	INVX1 X807 (.VDD(), .GND(), .A(G32), .Y());
	INVX1 X808 (.VDD(VDD), .GND(GND), .A(U486/a_13_43#), .Y(U486/a_18_54#));
	INVX1 X809 (.VDD(), .GND(), .A(G32), .Y());
	INVX1 X810 (.VDD(), .GND(), .A(U486/a_2_6#), .Y());
	INVX1 X811 (.VDD(), .GND(), .A(G28), .Y());
	INVX1 X812 (.VDD(VDD), .GND(GND), .A(G28), .Y(U486/a_13_43#));
	INVX1 X813 (.VDD(), .GND(), .A(n426), .Y());
	INVX1 X814 (.VDD(VDD), .GND(GND), .A(U487/a_13_43#), .Y(U487/a_18_54#));
	INVX1 X815 (.VDD(), .GND(), .A(n426), .Y());
	INVX1 X816 (.VDD(), .GND(), .A(U487/a_2_6#), .Y());
	INVX1 X817 (.VDD(), .GND(), .A(n421), .Y());
	INVX1 X818 (.VDD(VDD), .GND(GND), .A(n421), .Y(U487/a_13_43#));
	INVX1 X819 (.VDD(), .GND(), .A(n427), .Y());
	INVX1 X820 (.VDD(VDD), .GND(GND), .A(U488/a_12_41#), .Y(U488/a_18_54#));
	INVX1 X821 (.VDD(), .GND(), .A(U488/a_2_6#), .Y());
	INVX1 X822 (.VDD(), .GND(), .A(n427), .Y());
	INVX1 X823 (.VDD(), .GND(), .A(n428), .Y());
	INVX1 X824 (.VDD(VDD), .GND(GND), .A(n428), .Y(U488/a_12_41#));
	INVX1 X825 (.VDD(), .GND(), .A(G8), .Y());
	INVX1 X826 (.VDD(VDD), .GND(GND), .A(U489/a_13_43#), .Y(U489/a_18_54#));
	INVX1 X827 (.VDD(), .GND(), .A(G8), .Y());
	INVX1 X828 (.VDD(), .GND(), .A(U489/a_2_6#), .Y());
	INVX1 X829 (.VDD(), .GND(), .A(G7), .Y());
	INVX1 X830 (.VDD(VDD), .GND(GND), .A(G7), .Y(U489/a_13_43#));
	INVX1 X831 (.VDD(), .GND(), .A(G5), .Y());
	INVX1 X832 (.VDD(VDD), .GND(GND), .A(U490/a_12_41#), .Y(U490/a_18_54#));
	INVX1 X833 (.VDD(), .GND(), .A(U490/a_2_6#), .Y());
	INVX1 X834 (.VDD(), .GND(), .A(G5), .Y());
	INVX1 X835 (.VDD(), .GND(), .A(G6), .Y());
	INVX1 X836 (.VDD(VDD), .GND(GND), .A(G6), .Y(U490/a_12_41#));
	INVX1 X837 (.VDD(), .GND(), .A(n245), .Y());
	INVX1 X838 (.VDD(VDD), .GND(GND), .A(U491/a_13_43#), .Y(U491/a_18_54#));
	INVX1 X839 (.VDD(), .GND(), .A(n245), .Y());
	INVX1 X840 (.VDD(), .GND(), .A(U491/a_2_6#), .Y());
	INVX1 X841 (.VDD(), .GND(), .A(n430), .Y());
	INVX1 X842 (.VDD(VDD), .GND(GND), .A(n430), .Y(U491/a_13_43#));
	INVX1 X843 (.VDD(VDD), .GND(GND), .A(n290), .Y(n330));
	INVX1 X844 (.VDD(), .GND(), .A(n431), .Y());
	INVX1 X845 (.VDD(VDD), .GND(GND), .A(U493/a_12_41#), .Y(U493/a_18_54#));
	INVX1 X846 (.VDD(), .GND(), .A(U493/a_2_6#), .Y());
	INVX1 X847 (.VDD(), .GND(), .A(n431), .Y());
	INVX1 X848 (.VDD(), .GND(), .A(n432), .Y());
	INVX1 X849 (.VDD(VDD), .GND(GND), .A(n432), .Y(U493/a_12_41#));
	INVX1 X850 (.VDD(), .GND(), .A(n433), .Y());
	INVX1 X851 (.VDD(VDD), .GND(GND), .A(U494/a_13_43#), .Y(U494/a_18_54#));
	INVX1 X852 (.VDD(), .GND(), .A(n433), .Y());
	INVX1 X853 (.VDD(), .GND(), .A(U494/a_2_6#), .Y());
	INVX1 X854 (.VDD(), .GND(), .A(n434), .Y());
	INVX1 X855 (.VDD(VDD), .GND(GND), .A(n434), .Y(U494/a_13_43#));
	INVX1 X856 (.VDD(), .GND(), .A(G22), .Y());
	INVX1 X857 (.VDD(VDD), .GND(GND), .A(U495/a_13_43#), .Y(U495/a_18_54#));
	INVX1 X858 (.VDD(), .GND(), .A(G22), .Y());
	INVX1 X859 (.VDD(), .GND(), .A(U495/a_2_6#), .Y());
	INVX1 X860 (.VDD(), .GND(), .A(G18), .Y());
	INVX1 X861 (.VDD(VDD), .GND(GND), .A(G18), .Y(U495/a_13_43#));
	INVX1 X862 (.VDD(), .GND(), .A(G30), .Y());
	INVX1 X863 (.VDD(VDD), .GND(GND), .A(U496/a_13_43#), .Y(U496/a_18_54#));
	INVX1 X864 (.VDD(), .GND(), .A(G30), .Y());
	INVX1 X865 (.VDD(), .GND(), .A(U496/a_2_6#), .Y());
	INVX1 X866 (.VDD(), .GND(), .A(G26), .Y());
	INVX1 X867 (.VDD(VDD), .GND(GND), .A(G26), .Y(U496/a_13_43#));
	INVX1 X868 (.VDD(), .GND(), .A(n435), .Y());
	INVX1 X869 (.VDD(VDD), .GND(GND), .A(U497/a_13_43#), .Y(U497/a_18_54#));
	INVX1 X870 (.VDD(), .GND(), .A(n435), .Y());
	INVX1 X871 (.VDD(), .GND(), .A(U497/a_2_6#), .Y());
	INVX1 X872 (.VDD(), .GND(), .A(n374), .Y());
	INVX1 X873 (.VDD(VDD), .GND(GND), .A(n374), .Y(U497/a_13_43#));
	INVX1 X874 (.VDD(), .GND(), .A(n436), .Y());
	INVX1 X875 (.VDD(VDD), .GND(GND), .A(U498/a_12_41#), .Y(U498/a_18_54#));
	INVX1 X876 (.VDD(), .GND(), .A(U498/a_2_6#), .Y());
	INVX1 X877 (.VDD(), .GND(), .A(n436), .Y());
	INVX1 X878 (.VDD(), .GND(), .A(n437), .Y());
	INVX1 X879 (.VDD(VDD), .GND(GND), .A(n437), .Y(U498/a_12_41#));
	INVX1 X880 (.VDD(), .GND(), .A(G9), .Y());
	INVX1 X881 (.VDD(VDD), .GND(GND), .A(U499/a_13_43#), .Y(U499/a_18_54#));
	INVX1 X882 (.VDD(), .GND(), .A(G9), .Y());
	INVX1 X883 (.VDD(), .GND(), .A(U499/a_2_6#), .Y());
	INVX1 X884 (.VDD(), .GND(), .A(G12), .Y());
	INVX1 X885 (.VDD(VDD), .GND(GND), .A(G12), .Y(U499/a_13_43#));
	INVX1 X886 (.VDD(), .GND(), .A(G10), .Y());
	INVX1 X887 (.VDD(VDD), .GND(GND), .A(U500/a_12_41#), .Y(U500/a_18_54#));
	INVX1 X888 (.VDD(), .GND(), .A(U500/a_2_6#), .Y());
	INVX1 X889 (.VDD(), .GND(), .A(G10), .Y());
	INVX1 X890 (.VDD(), .GND(), .A(G11), .Y());
	INVX1 X891 (.VDD(VDD), .GND(GND), .A(G11), .Y(U500/a_12_41#));
	INVX1 X892 (.VDD(), .GND(), .A(n243), .Y());
	INVX1 X893 (.VDD(VDD), .GND(GND), .A(U501/a_13_43#), .Y(U501/a_18_54#));
	INVX1 X894 (.VDD(), .GND(), .A(n243), .Y());
	INVX1 X895 (.VDD(), .GND(), .A(U501/a_2_6#), .Y());
	INVX1 X896 (.VDD(), .GND(), .A(n430), .Y());
	INVX1 X897 (.VDD(VDD), .GND(GND), .A(n430), .Y(U501/a_13_43#));
	INVX1 X898 (.VDD(), .GND(), .A(n439), .Y());
	INVX1 X899 (.VDD(VDD), .GND(GND), .A(U502/a_12_41#), .Y(U502/a_18_54#));
	INVX1 X900 (.VDD(), .GND(), .A(U502/a_2_6#), .Y());
	INVX1 X901 (.VDD(), .GND(), .A(n439), .Y());
	INVX1 X902 (.VDD(), .GND(), .A(n440), .Y());
	INVX1 X903 (.VDD(VDD), .GND(GND), .A(n440), .Y(U502/a_12_41#));
	INVX1 X904 (.VDD(), .GND(), .A(G16), .Y());
	INVX1 X905 (.VDD(VDD), .GND(GND), .A(U503/a_13_43#), .Y(U503/a_18_54#));
	INVX1 X906 (.VDD(), .GND(), .A(G16), .Y());
	INVX1 X907 (.VDD(), .GND(), .A(U503/a_2_6#), .Y());
	INVX1 X908 (.VDD(), .GND(), .A(G15), .Y());
	INVX1 X909 (.VDD(VDD), .GND(GND), .A(G15), .Y(U503/a_13_43#));
	INVX1 X910 (.VDD(), .GND(), .A(G13), .Y());
	INVX1 X911 (.VDD(VDD), .GND(GND), .A(U504/a_12_41#), .Y(U504/a_18_54#));
	INVX1 X912 (.VDD(), .GND(), .A(U504/a_2_6#), .Y());
	INVX1 X913 (.VDD(), .GND(), .A(G13), .Y());
	INVX1 X914 (.VDD(), .GND(), .A(G14), .Y());
	INVX1 X915 (.VDD(VDD), .GND(GND), .A(G14), .Y(U504/a_12_41#));
endmodule
