module c1(inout A, inout AN, inout VDD, inout GND)
	INVERTER X1 (.A(A), .AN(AN), .VDD(VDD), .GND());
endmodule
