module c1355(inout G1, inout G10, inout G11, inout G12, inout G13, inout N384, inout N385, inout N386, inout N387, inout N388, inout N389, inout N390, inout N391, inout N392, inout N393, inout N394, inout N395, inout N396, inout N397, inout N398, inout N399, inout N400, inout N401, inout N402, inout N403, inout N404, inout N405, inout N406, inout N407, inout N408, inout N409, inout N410, inout N411, inout N412, inout N413, inout N414, inout N415, inout G14, inout G15, inout G16, inout G17, inout G18, inout G19, inout G2, inout G20, inout G21, inout G22, inout G23, inout G24, inout G25, inout G26, inout G27, inout G28, inout G29, inout G3, inout G30, inout G31, inout G32, inout G33, inout G34, inout G35, inout G36, inout G37, inout G38, inout G39, inout G4, inout G40, inout G41, inout G5, inout G6, inout G7, inout G8, inout G9, inout VDD, inout GND)
	XNOR2X1 X1 (.A(n232), .B(n232), .Y(U254/a_2_6#), .VDD(VDD), .GND());
	XNOR2X1 X2 (.A(n231), .B(n233), .Y(n350), .VDD(U255/a_2_6#), .GND());
	XNOR2X1 X3 (.A(n293), .B(n304), .Y(GND), .VDD(VDD), .GND());
	XNOR2X1 X4 (.A(n304), .B(n314), .Y(VDD), .VDD(GND), .GND());
	XNOR2X1 X5 (.A(U259/a_2_6#), .B(U260/a_2_6#), .Y(n225), .VDD(n225), .GND());
	XNOR2X1 X6 (.A(U260/a_2_6#), .B(U261/a_2_6#), .Y(n227), .VDD(n226), .GND());
	XNOR2X1 X7 (.A(U262/a_2_6#), .B(U263/a_2_6#), .Y(n228), .VDD(n228), .GND());
	XNOR2X1 X8 (.A(U263/a_2_6#), .B(U264/a_2_6#), .Y(n230), .VDD(n229), .GND());
	XNOR2X1 X9 (.A(n375), .B(U266/a_2_6#), .Y(n232), .VDD(GND), .GND());
	XNOR2X1 X10 (.A(n376), .B(n307), .Y(VDD), .VDD(GND), .GND());
	XNOR2X1 X11 (.A(n306), .B(n316), .Y(VDD), .VDD(n234), .GND());
	XNOR2X1 X12 (.A(n315), .B(n286), .Y(VDD), .VDD(n235), .GND());
	XNOR2X1 X13 (.A(n351), .B(U282/a_2_6#), .Y(GND), .VDD(n236), .GND());
	XNOR2X1 X14 (.A(U274/a_2_54#), .B(n359), .Y(n359), .VDD(n359), .GND());
	XNOR2X1 X15 (.A(n350), .B(n353), .Y(VDD), .VDD(n239), .GND());
	XNOR2X1 X16 (.A(n356), .B(n344), .Y(VDD), .VDD(n240), .GND());
	XNOR2X1 X17 (.A(n346), .B(G36), .Y(VDD), .VDD(n241), .GND());
	XNOR2X1 X18 (.A(n391), .B(U284/a_2_6#), .Y(n438), .VDD(n242), .GND());
	XNOR2X1 X19 (.A(n438), .B(U286/a_2_6#), .Y(n420), .VDD(n243), .GND());
	XNOR2X1 X20 (.A(n420), .B(U288/a_2_6#), .Y(n429), .VDD(n244), .GND());
	XNOR2X1 X21 (.A(n429), .B(n362), .Y(GND), .VDD(n245), .GND());
	XNOR2X1 X22 (.A(n288), .B(n319), .Y(U292/a_2_6#), .VDD(VDD), .GND());
	XNOR2X1 X23 (.A(n320), .B(G41), .Y(VDD), .VDD(n247), .GND());
	XNOR2X1 X24 (.A(n373), .B(G35), .Y(VDD), .VDD(n248), .GND());
	XNOR2X1 X25 (.A(n410), .B(n361), .Y(VDD), .VDD(n249), .GND());
	XNOR2X1 X26 (.A(n360), .B(n353), .Y(VDD), .VDD(n250), .GND());
	XNOR2X1 X27 (.A(n355), .B(n344), .Y(VDD), .VDD(n251), .GND());
	XNOR2X1 X28 (.A(n340), .B(G7), .Y(n252), .VDD(GND), .GND());
	XNOR2X1 X29 (.A(n348), .B(U304/a_2_6#), .Y(n318), .VDD(n252), .GND());
	XNOR2X1 X30 (.A(n318), .B(n312), .Y(GND), .VDD(n253), .GND());
	XNOR2X1 X31 (.A(n292), .B(n300), .Y(U308/a_2_6#), .VDD(VDD), .GND());
	XNOR2X1 X32 (.A(n303), .B(n340), .Y(U310/a_2_6#), .VDD(n255), .GND());
	XNOR2X1 X33 (.A(n338), .B(U312/a_2_6#), .Y(U312/a_2_6#), .VDD(n256), .GND());
	XNOR2X1 X34 (.A(G41), .B(n353), .Y(n257), .VDD(GND), .GND());
	XNOR2X1 X35 (.A(U314/a_2_6#), .B(n352), .Y(GND), .VDD(n352), .GND());
	XNOR2X1 X36 (.A(n344), .B(n345), .Y(GND), .VDD(U316/a_2_6#), .GND());
	XNOR2X1 X37 (.A(n319), .B(n321), .Y(GND), .VDD(U318/a_2_6#), .GND());
	XNOR2X1 X38 (.A(U320/a_2_6#), .B(n300), .Y(GND), .VDD(n309), .GND());
	XNOR2X1 X39 (.A(U322/a_2_6#), .B(n285), .Y(n262), .VDD(n301), .GND());
	XNOR2X1 X40 (.A(n292), .B(U326/a_2_6#), .Y(U326/a_2_6#), .VDD(GND), .GND());
	XNOR2X1 X41 (.A(n400), .B(n336), .Y(U328/a_2_6#), .VDD(n264), .GND());
	XNOR2X1 X42 (.A(n354), .B(n307), .Y(n343), .VDD(n265), .GND());
	XNOR2X1 X43 (.A(n334), .B(n337), .Y(GND), .VDD(U332/a_2_6#), .GND());
	XNOR2X1 X44 (.A(U334/a_2_6#), .B(n310), .Y(GND), .VDD(n322), .GND());
	XNOR2X1 X45 (.A(U336/a_2_6#), .B(n300), .Y(n269), .VDD(n311), .GND());
	XNOR2X1 X46 (.A(n286), .B(n290), .Y(n270), .VDD(GND), .GND());
	XNOR2X1 X47 (.A(n361), .B(n364), .Y(n364), .VDD(U342/a_2_6#), .GND());
	XNOR2X1 X48 (.A(n334), .B(n307), .Y(n333), .VDD(U344/a_2_6#), .GND());
	XNOR2X1 X49 (.A(n333), .B(U346/a_2_6#), .Y(U346/a_2_6#), .VDD(n273), .GND());
	XNOR2X1 X50 (.A(n292), .B(U348/a_2_6#), .Y(U348/a_2_6#), .VDD(GND), .GND());
	XNOR2X1 X51 (.A(n286), .B(U350/a_2_6#), .Y(U350/a_2_6#), .VDD(GND), .GND());
	XNOR2X1 X52 (.A(n308), .B(n288), .Y(U352/a_2_6#), .VDD(n276), .GND());
	XNOR2X1 X53 (.A(n328), .B(n363), .Y(n363), .VDD(n277), .GND());
	XNOR2X1 X54 (.A(n334), .B(n290), .Y(n335), .VDD(VDD), .GND());
	XNOR2X1 X55 (.A(n300), .B(n302), .Y(n302), .VDD(n280), .GND());
	XNOR2X1 X56 (.A(n288), .B(U360/a_2_6#), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X57 (.A(n287), .B(n317), .Y(), .VDD(n281), .GND());
	XNOR2X1 X58 (.A(n286), .B(U364/a_2_6#), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X59 (.A(n331), .B(U366/a_2_6#), .Y(U366/a_18_54#), .VDD(n283), .GND());
	XNOR2X1 X60 (.A(G32), .B(n275), .Y(U366/a_18_6#), .VDD(U366/a_13_43#), .GND());
	XNOR2X1 X61 (.A(G32), .B(G31), .Y(), .VDD(U366/a_13_43#), .GND());
	XNOR2X1 X62 (.A(U367/a_13_43#), .B(G31), .Y(), .VDD(U367/a_18_6#), .GND());
	XNOR2X1 X63 (.A(U368/a_13_43#), .B(G30), .Y(), .VDD(U368/a_18_54#), .GND());
	XNOR2X1 X64 (.A(U368/a_13_43#), .B(G30), .Y(), .VDD(U368/a_18_6#), .GND());
	XNOR2X1 X65 (.A(U369/a_13_43#), .B(G29), .Y(), .VDD(U369/a_18_54#), .GND());
	XNOR2X1 X66 (.A(U369/a_13_43#), .B(G29), .Y(), .VDD(U369/a_18_6#), .GND());
	XNOR2X1 X67 (.A(n222), .B(n294), .Y(VDD), .VDD(n285), .GND());
	XNOR2X1 X68 (.A(n296), .B(n298), .Y(), .VDD(n296), .GND());
	XNOR2X1 X69 (.A(U373/a_2_6#), .B(U373/a_13_43#), .Y(U373/a_13_43#), .VDD(U373/a_18_6#), .GND());
	XNOR2X1 X70 (.A(n270), .B(U374/a_13_43#), .Y(U373/a_13_43#), .VDD(U374/a_18_54#), .GND());
	XNOR2X1 X71 (.A(U374/a_2_6#), .B(U374/a_13_43#), .Y(U374/a_13_43#), .VDD(U374/a_18_6#), .GND());
	XNOR2X1 X72 (.A(G27), .B(G26), .Y(U375/a_18_54#), .VDD(U374/a_13_43#), .GND());
	XNOR2X1 X73 (.A(U375/a_13_43#), .B(U376/a_13_43#), .Y(U375/a_13_43#), .VDD(U375/a_18_6#), .GND());
	XNOR2X1 X74 (.A(G25), .B(n255), .Y(U376/a_18_6#), .VDD(U376/a_13_43#), .GND());
	XNOR2X1 X75 (.A(G25), .B(n238), .Y(n300), .VDD(U376/a_13_43#), .GND());
	XNOR2X1 X76 (.A(n295), .B(U379/a_2_6#), .Y(), .VDD(U378/a_9_6#), .GND());
	XNOR2X1 X77 (.A(G24), .B(G24), .Y(), .VDD(U379/a_13_43#), .GND());
	XNOR2X1 X78 (.A(U380/a_2_6#), .B(U380/a_13_43#), .Y(U380/a_13_43#), .VDD(U380/a_18_6#), .GND());
	XNOR2X1 X79 (.A(n269), .B(U381/a_13_43#), .Y(U380/a_13_43#), .VDD(U381/a_18_54#), .GND());
	XNOR2X1 X80 (.A(U381/a_2_6#), .B(n254), .Y(U381/a_13_43#), .VDD(), .GND());
	XNOR2X1 X81 (.A(G22), .B(G21), .Y(), .VDD(U381/a_13_43#), .GND());
	XNOR2X1 X82 (.A(n274), .B(n224), .Y(U382/a_13_43#), .VDD(n310), .GND());
	XNOR2X1 X83 (.A(n238), .B(U385/a_13_43#), .Y(U384/a_9_6#), .VDD(VDD), .GND());
	XNOR2X1 X84 (.A(U385/a_2_6#), .B(n253), .Y(U385/a_13_43#), .VDD(), .GND());
	XNOR2X1 X85 (.A(G20), .B(G19), .Y(), .VDD(U385/a_13_43#), .GND());
	XNOR2X1 X86 (.A(n247), .B(U387/a_13_43#), .Y(U386/a_13_43#), .VDD(U387/a_18_54#), .GND());
	XNOR2X1 X87 (.A(U387/a_2_6#), .B(n260), .Y(U387/a_13_43#), .VDD(), .GND());
	XNOR2X1 X88 (.A(G18), .B(U388/a_2_6#), .Y(U388/a_18_54#), .VDD(U387/a_13_43#), .GND());
	XNOR2X1 X89 (.A(G17), .B(n268), .Y(U388/a_18_6#), .VDD(U388/a_13_43#), .GND());
	XNOR2X1 X90 (.A(G17), .B(n298), .Y(n319), .VDD(U388/a_13_43#), .GND());
	XNOR2X1 X91 (.A(n297), .B(n295), .Y(), .VDD(U390/a_9_6#), .GND());
	XNOR2X1 X92 (.A(n305), .B(n305), .Y(GND), .VDD(GND), .GND());
	XNOR2X1 X93 (.A(n327), .B(n277), .Y(n326), .VDD(n326), .GND());
	XNOR2X1 X94 (.A(n330), .B(n283), .Y(n325), .VDD(n325), .GND());
	XNOR2X1 X95 (.A(n273), .B(G16), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X96 (.A(n273), .B(G16), .Y(), .VDD(GND), .GND());
	XNOR2X1 X97 (.A(n279), .B(G15), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X98 (.A(n279), .B(G15), .Y(), .VDD(GND), .GND());
	XNOR2X1 X99 (.A(n267), .B(G14), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X100 (.A(n267), .B(G14), .Y(), .VDD(GND), .GND());
	XNOR2X1 X101 (.A(n256), .B(n339), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X102 (.A(n256), .B(n339), .Y(), .VDD(GND), .GND());
	XNOR2X1 X103 (.A(n226), .B(n332), .Y(n341), .VDD(n334), .GND());
	XNOR2X1 X104 (.A(n329), .B(n329), .Y(), .VDD(n342), .GND());
	XNOR2X1 X105 (.A(U401/a_13_43#), .B(G12), .Y(), .VDD(U401/a_18_54#), .GND());
	XNOR2X1 X106 (.A(U401/a_13_43#), .B(U402/a_13_43#), .Y(), .VDD(U401/a_18_6#), .GND());
	XNOR2X1 X107 (.A(U402/a_2_6#), .B(n259), .Y(U402/a_18_6#), .VDD(), .GND());
	XNOR2X1 X108 (.A(U403/a_12_41#), .B(n347), .Y(), .VDD(U403/a_18_54#), .GND());
	XNOR2X1 X109 (.A(U403/a_12_41#), .B(n347), .Y(), .VDD(U403/a_18_6#), .GND());
	XNOR2X1 X110 (.A(U404/a_13_43#), .B(U404/a_13_43#), .Y(), .VDD(U404/a_18_54#), .GND());
	XNOR2X1 X111 (.A(n252), .B(n227), .Y(U404/a_13_43#), .VDD(n344), .GND());
	XNOR2X1 X112 (.A(n239), .B(n236), .Y(U406/a_9_6#), .VDD(VDD), .GND());
	XNOR2X1 X113 (.A(U407/a_13_43#), .B(G8), .Y(), .VDD(U407/a_18_54#), .GND());
	XNOR2X1 X114 (.A(U407/a_13_43#), .B(G8), .Y(), .VDD(U407/a_18_6#), .GND());
	XNOR2X1 X115 (.A(U408/a_13_43#), .B(G7), .Y(), .VDD(U408/a_18_54#), .GND());
	XNOR2X1 X116 (.A(U408/a_2_6#), .B(n251), .Y(VDD), .VDD(), .GND());
	XNOR2X1 X117 (.A(n251), .B(G6), .Y(), .VDD(GND), .GND());
	XNOR2X1 X118 (.A(n240), .B(n240), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X119 (.A(n240), .B(n228), .Y(GND), .VDD(n353), .GND());
	XNOR2X1 X120 (.A(n330), .B(n239), .Y(n358), .VDD(n358), .GND());
	XNOR2X1 X121 (.A(n250), .B(G4), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X122 (.A(n250), .B(G4), .Y(), .VDD(GND), .GND());
	XNOR2X1 X123 (.A(n246), .B(G3), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X124 (.A(n246), .B(G3), .Y(), .VDD(GND), .GND());
	XNOR2X1 X125 (.A(n278), .B(G2), .Y(), .VDD(VDD), .GND());
	XNOR2X1 X126 (.A(n278), .B(G2), .Y(), .VDD(GND), .GND());
	NOR3X1 X127 (.VDD(VDD), .GND(), .A(n375), .B(G38), .C(), .Y());
	NOR3X1 X128 (.VDD(VDD), .GND(), .A(n326), .B(G41), .C(), .Y());
	NOR3X1 X129 (.VDD(), .GND(), .A(n282), .B(n361), .C(), .Y());
	NOR3X1 X130 (.VDD(), .GND(), .A(n286), .B(G37), .C(), .Y());
	NOR3X1 X131 (.VDD(U280/a_2_6#), .GND(), .A(n344), .B(G39), .C(), .Y());
	NOR3X1 X132 (.VDD(VDD), .GND(), .A(n316), .B(G35), .C(), .Y());
	NOR3X1 X133 (.VDD(U282/a_2_6#), .GND(), .A(G36), .B(n307), .C(), .Y());
	NOR3X1 X134 (.VDD(), .GND(), .A(G41), .B(n316), .C(), .Y());
	NOR3X1 X135 (.VDD(U373/a_18_54#), .GND(), .A(U373/a_13_43#), .B(U375/a_2_6#), .C(), .Y());
	NOR3X1 X136 (.VDD(), .GND(), .A(n255), .B(U379/a_13_43#), .C(), .Y());
	NOR3X1 X137 (.VDD(), .GND(), .A(n274), .B(U385/a_13_43#), .C(), .Y());
	NOR3X1 X138 (.VDD(U382/a_18_6#), .GND(), .A(U382/a_13_43#), .B(n253), .C(), .Y());
	NOR3X1 X139 (.VDD(), .GND(), .A(n247), .B(U387/a_13_43#), .C(), .Y());
	NOR3X1 X140 (.VDD(), .GND(), .A(n350), .B(G11), .C(), .Y());
	NOR3X1 X141 (.VDD(), .GND(), .A(n350), .B(G12), .C(), .Y());
	NOR3X1 X142 (.VDD(U409/a_13_43#), .GND(), .A(G6), .B(n357), .C(), .Y());
	NAND3X1 X143 (.VDD(n343), .GND(), .A(n292), .B(U330/a_2_6#), .C(n343), .Y(GND));
	NAND3X1 X144 (.VDD(U372/a_2_64#), .GND(), .A(n286), .B(n297), .C(n297), .Y(VDD));
	NAND3X1 X145 (.VDD(GND), .GND(), .A(n299), .B(n285), .C(U367/a_13_43#), .Y(n270));
	NAND3X1 X146 (.VDD(VDD), .GND(), .A(U340/a_2_6#), .B(n285), .C(n313), .Y(n289));
	NAND3X1 X147 (.VDD(GND), .GND(), .A(U354/a_2_6#), .B(n307), .C(U362/a_2_6#), .Y(n363));
	NAND3X1 X148 (.VDD(n341), .GND(), .A(n254), .B(n342), .C(n332), .Y(VDD));
	BUFX2 X149 (.VDD(n338), .GND(), .A(U310/a_2_6#), .Y());
	BUFX2 X150 (.VDD(n345), .GND(), .A(U316/a_2_6#), .Y());
	BUFX2 X151 (.VDD(VDD), .GND(), .A(n290), .Y(n321));
	BUFX2 X152 (.VDD(n260), .GND(), .A(n321), .Y(U320/a_2_6#));
	BUFX2 X153 (.VDD(n309), .GND(), .A(U320/a_2_6#), .Y(n261));
	BUFX2 X154 (.VDD(), .GND(), .A(n300), .Y());
	BUFX2 X155 (.VDD(n291), .GND(), .A(U324/a_2_6#), .Y(n263));
	BUFX2 X156 (.VDD(), .GND(), .A(G33), .Y());
	BUFX2 X157 (.VDD(VDD), .GND(), .A(n336), .Y(n354));
	BUFX2 X158 (.VDD(n265), .GND(), .A(n354), .Y(U330/a_2_6#));
	BUFX2 X159 (.VDD(VDD), .GND(), .A(n316), .Y(n337));
	BUFX2 X160 (.VDD(n267), .GND(), .A(n337), .Y(U334/a_2_6#));
	BUFX2 X161 (.VDD(n322), .GND(), .A(U334/a_2_6#), .Y(n268));
	BUFX2 X162 (.VDD(), .GND(), .A(n310), .Y());
	BUFX2 X163 (.VDD(n271), .GND(), .A(n289), .Y(n271));
	BUFX2 X164 (.VDD(GND), .GND(), .A(n340), .Y(n364));
	BUFX2 X165 (.VDD(n284), .GND(), .A(U348/a_2_6#), .Y(n275));
	BUFX2 X166 (.VDD(), .GND(), .A(n336), .Y());
	BUFX2 X167 (.VDD(VDD), .GND(), .A(n288), .Y(n328));
	BUFX2 X168 (.VDD(n277), .GND(), .A(n328), .Y(U354/a_2_6#));
	BUFX2 X169 (.VDD(VDD), .GND(), .A(n336), .Y(n335));
	BUFX2 X170 (.VDD(n279), .GND(), .A(n335), .Y(U358/a_2_6#));
	BUFX2 X171 (.VDD(n317), .GND(), .A(U362/a_2_6#), .Y(n282));
	BUFX2 X172 (.VDD(GND), .GND(), .A(n298), .Y(n296));
	BUFX2 X173 (.VDD(), .GND(), .A(U374/a_2_6#), .Y());
	BUFX2 X174 (.VDD(), .GND(), .A(U375/a_2_6#), .Y());
	BUFX2 X175 (.VDD(VDD), .GND(), .A(n261), .Y(U379/a_18_54#));
	BUFX2 X176 (.VDD(VDD), .GND(), .A(n269), .Y(U380/a_18_54#));
	BUFX2 X177 (.VDD(VDD), .GND(), .A(n247), .Y(U386/a_18_54#));
	BUFX2 X178 (.VDD(U402/a_13_43#), .GND(), .A(G11), .Y());
	BUFX2 X179 (.VDD(U404/a_13_43#), .GND(), .A(G9), .Y());
	INVX1 X180 (.VDD(), .GND(), .A(n230), .Y());
	INVX1 X181 (.VDD(), .GND(), .A(n376), .Y());
	INVX1 X182 (.VDD(), .GND(), .A(n307), .Y());
	INVX1 X183 (.VDD(), .GND(), .A(n276), .Y());
	INVX1 X184 (.VDD(), .GND(), .A(n316), .Y());
	INVX1 X185 (.VDD(), .GND(), .A(n288), .Y());
	INVX1 X186 (.VDD(), .GND(), .A(G41), .Y());
	INVX1 X187 (.VDD(VDD), .GND(), .A(n361), .Y(U290/a_2_6#));
	INVX1 X188 (.VDD(), .GND(), .A(n336), .Y());
	INVX1 X189 (.VDD(VDD), .GND(), .A(G41), .Y(U294/a_2_6#));
	INVX1 X190 (.VDD(VDD), .GND(), .A(n353), .Y(U300/a_2_6#));
	INVX1 X191 (.VDD(VDD), .GND(), .A(n344), .Y(U302/a_2_6#));
	INVX1 X192 (.VDD(VDD), .GND(), .A(n319), .Y(U304/a_2_6#));
	INVX1 X193 (.VDD(), .GND(), .A(n286), .Y());
	INVX1 X194 (.VDD(VDD), .GND(), .A(n310), .Y(U306/a_2_6#));
	INVX1 X195 (.VDD(), .GND(), .A(n290), .Y());
	INVX1 X196 (.VDD(), .GND(), .A(n292), .Y());
	INVX1 X197 (.VDD(VDD), .GND(), .A(U324/a_2_6#), .Y(n291));
	INVX1 X198 (.VDD(VDD), .GND(), .A(U338/a_2_6#), .Y(n299));
	INVX1 X199 (.VDD(GND), .GND(), .A(n313), .Y(n274));
	INVX1 X200 (.VDD(VDD), .GND(), .A(n363), .Y(n278));
	INVX1 X201 (.VDD(), .GND(), .A(n281), .Y());
	INVX1 X202 (.VDD(), .GND(), .A(n270), .Y());
	INVX1 X203 (.VDD(), .GND(), .A(U376/a_2_6#), .Y());
	INVX1 X204 (.VDD(GND), .GND(), .A(U381/a_13_43#), .Y(U381/a_18_6#));
	INVX1 X205 (.VDD(VDD), .GND(), .A(U382/a_13_43#), .Y(U382/a_18_54#));
	INVX1 X206 (.VDD(), .GND(), .A(n274), .Y());
	INVX1 X207 (.VDD(GND), .GND(), .A(U386/a_13_43#), .Y(U386/a_18_6#));
	INVX1 X208 (.VDD(VDD), .GND(), .A(n329), .Y(U400/a_2_64#));
	INVX1 X209 (.VDD(GND), .GND(), .A(n330), .Y(n342));
	INVX1 X210 (.VDD(), .GND(), .A(G6), .Y());
endmodule
