.SUBCKT c1355 G1 G10 G11 G12 G13 N384 N385 N386 N387 N388 N389 N390 N391 N392 N393 N394 N395 N396 N397 N398 N399 N400 N401 N402 N403 N404 N405 N406 N407 N408 N409 N410 N411 N412 N413 N414 N415 G14 G15 G16 G17 G18 G19 G2 G20 G21 G22 G23 G24 G25 G26 G27 G28 G29 G3 G30 G31 G32 G33 G34 G35 G36 G37 G38 G39 G4 G40 G41 G5 G6 G7 G8 G9 VDD GND 
M1 U254/a_2_6# n230 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M2 VDD n232 U254/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M3 n305 U254/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M4 U254/a_9_6# n230 U254/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M5 GND n232 U254/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M6 n305 U254/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M7 U255/a_2_6# n231 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M8 VDD n233 U255/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M9 n350 U255/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M10 U255/a_9_6# n231 U255/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M11 GND n233 U255/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M12 n350 U255/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M13 VDD n293 U256/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M14 n222 U256/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M15 GND n293 U256/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M16 n222 U256/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M17 VDD n304 U257/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M18 n223 U257/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M19 GND n304 U257/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M20 n223 U257/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M21 VDD n314 U258/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M22 n224 U258/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M23 GND n314 U258/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M24 n224 U258/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M25 VDD n323 U259/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M26 n225 U259/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M27 GND n323 U259/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M28 n225 U259/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M29 VDD n341 U260/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M30 n226 U260/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M31 GND n341 U260/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M32 n226 U260/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M33 VDD n349 U261/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M34 n227 U261/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M35 GND n349 U261/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M36 n227 U261/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M37 VDD n358 U262/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M38 n228 U262/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M39 GND n358 U262/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M40 n228 U262/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M41 VDD n365 U263/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M42 n229 U263/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M43 GND n365 U263/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M44 n229 U263/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M45 VDD n325 U264/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M46 n230 U264/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M47 GND n325 U264/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M48 n230 U264/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M49 VDD n375 U265/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M50 n231 U265/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M51 GND n375 U265/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M52 n231 U265/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M53 VDD n326 U266/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M54 n232 U266/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M55 GND n326 U266/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M56 n232 U266/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M57 VDD n376 U267/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M58 n233 U267/a_2_6# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M59 GND n376 U267/a_2_6# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M60 n233 U267/a_2_6# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M61 U268/a_9_54# n307 U268/a_2_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M62 VDD n276 U268/a_9_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M63 n306 U268/a_2_54# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M64 U268/a_2_54# n307 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M65 GND n276 U268/a_2_54# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M66 n306 U268/a_2_54# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M67 n234 n306 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M68 n234 n306 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M69 U270/a_9_54# n316 U270/a_2_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M70 VDD n282 U270/a_9_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M71 n315 U270/a_2_54# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M72 U270/a_2_54# n316 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M73 GND n282 U270/a_2_54# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M74 n315 U270/a_2_54# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M75 n235 n315 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M76 n235 n315 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M77 U272/a_9_54# n286 U272/a_2_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M78 VDD n277 U272/a_9_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M79 n351 U272/a_2_54# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M80 U272/a_2_54# n286 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M81 GND n277 U272/a_2_54# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M82 n351 U272/a_2_54# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M83 n236 n351 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M84 n236 n351 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M85 U274/a_9_54# n288 U274/a_2_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M86 VDD n283 U274/a_9_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M87 n359 U274/a_2_54# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M88 U274/a_2_54# n288 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M89 GND n283 U274/a_2_54# GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M90 n359 U274/a_2_54# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M91 n237 n359 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M92 n237 n359 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M93 n238 n305 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M94 n238 n305 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M95 n239 n350 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M96 n239 n350 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M97 U278/a_2_6# n353 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M98 VDD n340 U278/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M99 n356 U278/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M100 U278/a_9_6# n353 U278/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M101 GND n340 U278/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M102 n356 U278/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M103 n240 n356 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M104 n240 n356 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M105 U280/a_2_6# n344 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M106 VDD n316 U280/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M107 n346 U280/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M108 U280/a_9_6# n344 U280/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M109 GND n316 U280/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M110 n346 U280/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M111 n241 n346 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M112 n241 n346 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M113 U282/a_2_6# G36 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M114 VDD G41 U282/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M115 n391 U282/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M116 U282/a_9_6# G36 U282/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M117 GND G41 U282/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M118 n391 U282/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M119 n242 n391 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M120 n242 n391 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M121 U284/a_2_6# G38 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M122 VDD G41 U284/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M123 n438 U284/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M124 U284/a_9_6# G38 U284/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M125 GND G41 U284/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M126 n438 U284/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M127 n243 n438 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M128 n243 n438 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M129 U286/a_2_6# G37 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M130 VDD G41 U286/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M131 n420 U286/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M132 U286/a_9_6# G37 U286/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M133 GND G41 U286/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M134 n420 U286/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M135 n244 n420 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M136 n244 n420 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M137 U288/a_2_6# G40 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M138 VDD G41 U288/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M139 n429 U288/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M140 U288/a_9_6# G40 U288/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M141 GND G41 U288/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M142 n429 U288/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M143 n245 n429 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M144 n245 n429 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M145 U290/a_2_6# n361 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M146 VDD n336 U290/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M147 n362 U290/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M148 U290/a_9_6# n361 U290/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M149 GND n336 U290/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M150 n362 U290/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M151 n246 n362 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M152 n246 n362 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M153 U292/a_2_6# n319 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M154 VDD n288 U292/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M155 n320 U292/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M156 U292/a_9_6# n319 U292/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M157 GND n288 U292/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M158 n320 U292/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M159 n247 n320 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M160 n247 n320 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M161 U294/a_2_6# G41 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M162 VDD G39 U294/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M163 n373 U294/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M164 U294/a_9_6# G41 U294/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M165 GND G39 U294/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M166 n373 U294/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M167 n248 n373 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M168 n248 n373 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M169 U296/a_2_6# G35 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M170 VDD G41 U296/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M171 n410 U296/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M172 U296/a_9_6# G35 U296/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M173 GND G41 U296/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M174 n410 U296/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M175 n249 n410 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M176 n249 n410 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M177 U298/a_2_6# n361 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M178 VDD n307 U298/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M179 n360 U298/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M180 U298/a_9_6# n361 U298/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M181 GND n307 U298/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M182 n360 U298/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M183 n250 n360 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M184 n250 n360 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M185 U300/a_2_6# n353 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M186 VDD n316 U300/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M187 n355 U300/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M188 U300/a_9_6# n353 U300/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M189 GND n316 U300/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M190 n355 U300/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M191 n251 n355 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M192 n251 n355 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M193 U302/a_2_6# n344 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M194 VDD n340 U302/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M195 n348 U302/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M196 U302/a_9_6# n344 U302/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M197 GND n340 U302/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M198 n348 U302/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M199 n252 n348 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M200 n252 n348 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M201 U304/a_2_6# n319 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M202 VDD n286 U304/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M203 n318 U304/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M204 U304/a_9_6# n319 U304/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M205 GND n286 U304/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M206 n318 U304/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M207 n253 n318 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M208 n253 n318 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M209 U306/a_2_6# n310 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M210 VDD n290 U306/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M211 n312 U306/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M212 U306/a_9_6# n310 U306/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M213 GND n290 U306/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M214 n312 U306/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M215 n254 n312 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M216 n254 n312 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M217 U308/a_2_6# n300 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M218 VDD n292 U308/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M219 n303 U308/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M220 U308/a_9_6# n300 U308/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M221 GND n292 U308/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M222 n303 U308/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M223 n255 n303 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M224 n255 n303 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M225 U310/a_2_6# n334 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M226 VDD n340 U310/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M227 n338 U310/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M228 U310/a_9_6# n334 U310/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M229 GND n340 U310/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M230 n338 U310/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M231 n256 n338 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M232 n256 n338 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M233 U312/a_2_6# G34 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M234 VDD G41 U312/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M235 n383 U312/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M236 U312/a_9_6# G34 U312/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M237 GND G41 U312/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M238 n383 U312/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M239 n257 n383 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M240 n257 n383 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M241 U314/a_2_6# n353 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M242 VDD n307 U314/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M243 n352 U314/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M244 U314/a_9_6# n353 U314/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M245 GND n307 U314/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M246 n352 U314/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M247 n258 n352 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M248 n258 n352 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M249 U316/a_2_6# n344 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M250 VDD n336 U316/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M251 n345 U316/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M252 U316/a_9_6# n344 U316/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M253 GND n336 U316/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M254 n345 U316/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M255 n259 n345 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M256 n259 n345 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M257 U318/a_2_6# n319 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M258 VDD n290 U318/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M259 n321 U318/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M260 U318/a_9_6# n319 U318/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M261 GND n290 U318/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M262 n321 U318/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M263 n260 n321 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M264 n260 n321 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M265 U320/a_2_6# n310 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M266 VDD n286 U320/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M267 n309 U320/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M268 U320/a_9_6# n310 U320/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M269 GND n286 U320/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M270 n309 U320/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M271 n261 n309 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M272 n261 n309 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M273 U322/a_2_6# n300 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M274 VDD n288 U322/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M275 n301 U322/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M276 U322/a_9_6# n300 U322/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M277 GND n288 U322/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M278 n301 U322/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M279 n262 n301 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M280 n262 n301 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M281 U324/a_2_6# n285 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M282 VDD n292 U324/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M283 n291 U324/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M284 U324/a_9_6# n285 U324/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M285 GND n292 U324/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M286 n291 U324/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M287 n263 n291 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M288 n263 n291 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M289 U326/a_2_6# G33 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M290 VDD G41 U326/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M291 n400 U326/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M292 U326/a_9_6# G33 U326/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M293 GND G41 U326/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M294 n400 U326/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M295 n264 n400 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M296 n264 n400 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M297 U328/a_2_6# n353 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M298 VDD n336 U328/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M299 n354 U328/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M300 U328/a_9_6# n353 U328/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M301 GND n336 U328/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M302 n354 U328/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M303 n265 n354 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M304 n265 n354 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M305 U330/a_2_6# n344 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M306 VDD n307 U330/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M307 n343 U330/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M308 U330/a_9_6# n344 U330/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M309 GND n307 U330/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M310 n343 U330/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M311 n266 n343 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M312 n266 n343 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M313 U332/a_2_6# n334 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M314 VDD n316 U332/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M315 n337 U332/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M316 U332/a_9_6# n334 U332/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M317 GND n316 U332/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M318 n337 U332/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M319 n267 n337 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M320 n267 n337 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M321 U334/a_2_6# n319 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M322 VDD n292 U334/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M323 n322 U334/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M324 U334/a_9_6# n319 U334/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M325 GND n292 U334/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M326 n322 U334/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M327 n268 n322 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M328 n268 n322 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M329 U336/a_2_6# n310 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M330 VDD n288 U336/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M331 n311 U336/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M332 U336/a_9_6# n310 U336/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M333 GND n288 U336/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M334 n311 U336/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M335 n269 n311 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M336 n269 n311 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M337 U338/a_2_6# n300 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M338 VDD n286 U338/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M339 n299 U338/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M340 U338/a_9_6# n300 U338/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M341 GND n286 U338/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M342 n299 U338/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M343 n270 n299 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M344 n270 n299 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M345 U340/a_2_6# n285 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M346 VDD n290 U340/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M347 n289 U340/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M348 U340/a_9_6# n285 U340/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M349 GND n290 U340/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M350 n289 U340/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M351 n271 n289 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M352 n271 n289 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M353 U342/a_2_6# n361 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M354 VDD n340 U342/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M355 n364 U342/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M356 U342/a_9_6# n361 U342/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M357 GND n340 U342/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M358 n364 U342/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M359 n272 n364 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M360 n272 n364 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M361 U344/a_2_6# n334 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M362 VDD n307 U344/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M363 n333 U344/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M364 U344/a_9_6# n334 U344/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M365 GND n307 U344/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M366 n333 U344/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M367 n273 n333 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M368 n273 n333 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M369 U346/a_2_6# n310 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M370 VDD n292 U346/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M371 n313 U346/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M372 U346/a_9_6# n310 U346/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M373 GND n292 U346/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M374 n313 U346/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M375 n274 n313 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M376 n274 n313 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M377 U348/a_2_6# n285 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M378 VDD n286 U348/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M379 n284 U348/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M380 U348/a_9_6# n285 U348/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M381 GND n286 U348/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M382 n284 U348/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M383 n275 n284 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M384 n275 n284 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M385 U350/a_2_6# n336 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M386 VDD n316 U350/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M387 n308 U350/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M388 U350/a_9_6# n336 U350/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M389 GND n316 U350/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M390 n308 U350/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M391 n276 n308 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M392 n276 n308 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M393 U352/a_2_6# n290 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M394 VDD n288 U352/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M395 n328 U352/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M396 U352/a_9_6# n290 U352/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M397 GND n288 U352/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M398 n328 U352/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M399 n277 n328 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M400 n277 n328 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M401 U354/a_2_6# n361 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M402 VDD n316 U354/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M403 n363 U354/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M404 U354/a_9_6# n361 U354/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M405 GND n316 U354/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M406 n363 U354/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M407 n278 n363 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M408 n278 n363 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M409 U356/a_2_6# n334 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M410 VDD n336 U356/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M411 n335 U356/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M412 U356/a_9_6# n334 U356/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M413 GND n336 U356/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M414 n335 U356/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M415 n279 n335 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M416 n279 n335 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M417 U358/a_2_6# n300 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M418 VDD n290 U358/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M419 n302 U358/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M420 U358/a_9_6# n300 U358/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M421 GND n290 U358/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M422 n302 U358/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M423 n280 n302 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M424 n280 n302 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M425 U360/a_2_6# n285 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M426 VDD n288 U360/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M427 n287 U360/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M428 U360/a_9_6# n285 U360/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M429 GND n288 U360/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M430 n287 U360/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M431 n281 n287 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M432 n281 n287 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M433 U362/a_2_6# n340 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M434 VDD n307 U362/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M435 n317 U362/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M436 U362/a_9_6# n340 U362/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M437 GND n307 U362/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M438 n317 U362/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M439 n282 n317 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M440 n282 n317 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M441 U364/a_2_6# n292 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M442 VDD n286 U364/a_2_6# VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M443 n331 U364/a_2_6# VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M444 U364/a_9_6# n292 U364/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M445 GND n286 U364/a_9_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M446 n331 U364/a_2_6# GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M447 n283 n331 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M448 n283 n331 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M449 VDD n275 U366/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M450 U366/a_18_54# U366/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M451 N415 n275 U366/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M452 U366/a_35_54# U366/a_2_6# N415 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M453 VDD G32 U366/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M454 U366/a_13_43# G32 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M455 GND n275 U366/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M456 U366/a_18_6# U366/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M457 N415 U366/a_2_6# U366/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M458 U366/a_35_6# n275 N415 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M459 GND G32 U366/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M460 U366/a_13_43# G32 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M461 VDD n281 U367/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M462 U367/a_18_54# U367/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M463 N414 n281 U367/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M464 U367/a_35_54# U367/a_2_6# N414 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M465 VDD G31 U367/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M466 U367/a_13_43# G31 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M467 GND n281 U367/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M468 U367/a_18_6# U367/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M469 N414 U367/a_2_6# U367/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M470 U367/a_35_6# n281 N414 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M471 GND G31 U367/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M472 U367/a_13_43# G31 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M473 VDD n271 U368/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M474 U368/a_18_54# U368/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M475 N413 n271 U368/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M476 U368/a_35_54# U368/a_2_6# N413 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M477 VDD G30 U368/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M478 U368/a_13_43# G30 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M479 GND n271 U368/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M480 U368/a_18_6# U368/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M481 N413 U368/a_2_6# U368/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M482 U368/a_35_6# n271 N413 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M483 GND G30 U368/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M484 U368/a_13_43# G30 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M485 VDD n263 U369/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M486 U369/a_18_54# U369/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M487 N412 n263 U369/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M488 U369/a_35_54# U369/a_2_6# N412 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M489 VDD G29 U369/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M490 U369/a_13_43# G29 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M491 GND n263 U369/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M492 U369/a_18_6# U369/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M493 N412 U369/a_2_6# U369/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M494 U369/a_35_6# n263 N412 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M495 GND G29 U369/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M496 U369/a_13_43# G29 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M497 n285 n222 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M498 n285 n222 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M499 n293 n294 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M500 VDD n295 n293 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M501 n293 n296 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M502 U371/a_9_6# n294 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M503 U371/a_14_6# n295 U371/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M504 n293 n296 U371/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M505 VDD n297 U372/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M506 U372/a_2_64# n297 VDD VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M507 U372/a_25_64# n305 U372/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M508 U372/a_2_64# n305 U372/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M509 n296 n298 U372/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M510 U372/a_25_64# n298 n296 VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M511 n296 n297 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M512 GND n305 n296 GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M513 n296 n298 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M514 VDD n270 U373/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M515 U373/a_18_54# U373/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M516 N411 n270 U373/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M517 U373/a_35_54# U373/a_2_6# N411 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M518 VDD G28 U373/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M519 U373/a_13_43# G28 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M520 GND n270 U373/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M521 U373/a_18_6# U373/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M522 N411 U373/a_2_6# U373/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M523 U373/a_35_6# n270 N411 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M524 GND G28 U373/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M525 U373/a_13_43# G28 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M526 VDD n262 U374/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M527 U374/a_18_54# U374/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M528 N410 n262 U374/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M529 U374/a_35_54# U374/a_2_6# N410 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M530 VDD G27 U374/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M531 U374/a_13_43# G27 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M532 GND n262 U374/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M533 U374/a_18_6# U374/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M534 N410 U374/a_2_6# U374/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M535 U374/a_35_6# n262 N410 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M536 GND G27 U374/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M537 U374/a_13_43# G27 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M538 VDD n280 U375/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M539 U375/a_18_54# U375/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M540 N409 n280 U375/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M541 U375/a_35_54# U375/a_2_6# N409 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M542 VDD G26 U375/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M543 U375/a_13_43# G26 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M544 GND n280 U375/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M545 U375/a_18_6# U375/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M546 N409 U375/a_2_6# U375/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M547 U375/a_35_6# n280 N409 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M548 GND G26 U375/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M549 U375/a_13_43# G26 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M550 VDD n255 U376/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M551 U376/a_18_54# U376/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M552 N408 n255 U376/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M553 U376/a_35_54# U376/a_2_6# N408 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M554 VDD G25 U376/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M555 U376/a_13_43# G25 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M556 GND n255 U376/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M557 U376/a_18_6# U376/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M558 N408 U376/a_2_6# U376/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M559 U376/a_35_6# n255 N408 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M560 GND G25 U376/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M561 U376/a_13_43# G25 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M562 n300 n223 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M563 n300 n223 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M564 n304 n295 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M565 VDD n238 n304 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M566 n304 n234 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M567 U378/a_9_6# n295 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M568 U378/a_14_6# n238 U378/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M569 n304 n234 U378/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M570 VDD n261 U379/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M571 U379/a_18_54# U379/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M572 N407 n261 U379/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M573 U379/a_35_54# U379/a_2_6# N407 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M574 VDD G24 U379/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M575 U379/a_13_43# G24 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M576 GND n261 U379/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M577 U379/a_18_6# U379/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M578 N407 U379/a_2_6# U379/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M579 U379/a_35_6# n261 N407 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M580 GND G24 U379/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M581 U379/a_13_43# G24 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M582 VDD n269 U380/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M583 U380/a_18_54# U380/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M584 N406 n269 U380/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M585 U380/a_35_54# U380/a_2_6# N406 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M586 VDD G23 U380/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M587 U380/a_13_43# G23 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M588 GND n269 U380/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M589 U380/a_18_6# U380/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M590 N406 U380/a_2_6# U380/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M591 U380/a_35_6# n269 N406 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M592 GND G23 U380/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M593 U380/a_13_43# G23 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M594 VDD n254 U381/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M595 U381/a_18_54# U381/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M596 N405 n254 U381/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M597 U381/a_35_54# U381/a_2_6# N405 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M598 VDD G22 U381/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M599 U381/a_13_43# G22 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M600 GND n254 U381/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M601 U381/a_18_6# U381/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M602 N405 U381/a_2_6# U381/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M603 U381/a_35_6# n254 N405 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M604 GND G22 U381/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M605 U381/a_13_43# G22 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M606 VDD n274 U382/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M607 U382/a_18_54# U382/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M608 N404 n274 U382/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M609 U382/a_35_54# U382/a_2_6# N404 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M610 VDD G21 U382/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M611 U382/a_13_43# G21 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M612 GND n274 U382/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M613 U382/a_18_6# U382/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M614 N404 U382/a_2_6# U382/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M615 U382/a_35_6# n274 N404 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M616 GND G21 U382/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M617 U382/a_13_43# G21 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M618 n310 n224 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M619 n310 n224 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M620 n314 n294 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M621 VDD n238 n314 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M622 n314 n235 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M623 U384/a_9_6# n294 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M624 U384/a_14_6# n238 U384/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M625 n314 n235 U384/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M626 VDD n253 U385/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M627 U385/a_18_54# U385/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M628 N403 n253 U385/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M629 U385/a_35_54# U385/a_2_6# N403 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M630 VDD G20 U385/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M631 U385/a_13_43# G20 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M632 GND n253 U385/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M633 U385/a_18_6# U385/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M634 N403 U385/a_2_6# U385/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M635 U385/a_35_6# n253 N403 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M636 GND G20 U385/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M637 U385/a_13_43# G20 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M638 VDD n247 U386/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M639 U386/a_18_54# U386/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M640 N402 n247 U386/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M641 U386/a_35_54# U386/a_2_6# N402 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M642 VDD G19 U386/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M643 U386/a_13_43# G19 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M644 GND n247 U386/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M645 U386/a_18_6# U386/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M646 N402 U386/a_2_6# U386/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M647 U386/a_35_6# n247 N402 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M648 GND G19 U386/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M649 U386/a_13_43# G19 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M650 VDD n260 U387/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M651 U387/a_18_54# U387/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M652 N401 n260 U387/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M653 U387/a_35_54# U387/a_2_6# N401 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M654 VDD G18 U387/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M655 U387/a_13_43# G18 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M656 GND n260 U387/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M657 U387/a_18_6# U387/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M658 N401 U387/a_2_6# U387/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M659 U387/a_35_6# n260 N401 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M660 GND G18 U387/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M661 U387/a_13_43# G18 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M662 VDD n268 U388/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M663 U388/a_18_54# U388/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M664 N400 n268 U388/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M665 U388/a_35_54# U388/a_2_6# N400 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M666 VDD G17 U388/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M667 U388/a_13_43# G17 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M668 GND n268 U388/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M669 U388/a_18_6# U388/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M670 N400 U388/a_2_6# U388/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M671 U388/a_35_6# n268 N400 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M672 GND G17 U388/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M673 U388/a_13_43# G17 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M674 n319 n225 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M675 n319 n225 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M676 n323 n297 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M677 VDD n298 n323 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M678 n323 n324 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M679 U390/a_9_6# n297 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M680 U390/a_14_6# n298 U390/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M681 n323 n324 U390/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M682 VDD n295 U391/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M683 U391/a_2_64# n295 VDD VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M684 U391/a_25_64# n305 U391/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M685 U391/a_2_64# n305 U391/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M686 n324 n294 U391/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M687 U391/a_25_64# n294 n324 VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M688 n324 n295 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M689 GND n305 n324 GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M690 n324 n294 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M691 n326 n327 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M692 VDD n277 n326 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M693 n326 n329 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M694 U392/a_9_6# n327 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M695 U392/a_14_6# n277 U392/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M696 n326 n329 U392/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M697 n325 n330 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M698 VDD n283 n325 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M699 n325 n332 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M700 U393/a_9_6# n330 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M701 U393/a_14_6# n283 U393/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M702 n325 n332 U393/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M703 VDD n273 U394/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M704 U394/a_18_54# U394/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M705 N399 n273 U394/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M706 U394/a_35_54# U394/a_2_6# N399 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M707 VDD G16 U394/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M708 U394/a_13_43# G16 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M709 GND n273 U394/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M710 U394/a_18_6# U394/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M711 N399 U394/a_2_6# U394/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M712 U394/a_35_6# n273 N399 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M713 GND G16 U394/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M714 U394/a_13_43# G16 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M715 VDD n279 U395/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M716 U395/a_18_54# U395/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M717 N398 n279 U395/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M718 U395/a_35_54# U395/a_2_6# N398 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M719 VDD G15 U395/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M720 U395/a_13_43# G15 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M721 GND n279 U395/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M722 U395/a_18_6# U395/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M723 N398 U395/a_2_6# U395/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M724 U395/a_35_6# n279 N398 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M725 GND G15 U395/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M726 U395/a_13_43# G15 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M727 VDD n267 U396/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M728 U396/a_18_54# U396/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M729 N397 n267 U396/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M730 U396/a_35_54# U396/a_2_6# N397 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M731 VDD G14 U396/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M732 U396/a_13_43# G14 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M733 GND n267 U396/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M734 U396/a_18_6# U396/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M735 N397 U396/a_2_6# U396/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M736 U396/a_35_6# n267 N397 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M737 GND G14 U396/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M738 U396/a_13_43# G14 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M739 VDD n256 U397/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M740 U397/a_18_54# U397/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M741 N396 U397/a_2_6# U397/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M742 U397/a_35_54# n256 N396 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M743 VDD n339 U397/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M744 U397/a_12_41# n339 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M745 GND n256 U397/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M746 U397/a_18_6# U397/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M747 N396 n256 U397/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M748 U397/a_35_6# U397/a_2_6# N396 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M749 GND n339 U397/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M750 U397/a_12_41# n339 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M751 n334 n226 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M752 n334 n226 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M753 n341 n327 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M754 VDD n332 n341 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M755 n341 n342 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M756 U399/a_9_6# n327 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M757 U399/a_14_6# n332 U399/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M758 n341 n342 U399/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M759 VDD n329 U400/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M760 U400/a_2_64# n329 VDD VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M761 U400/a_25_64# n350 U400/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M762 U400/a_2_64# n350 U400/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M763 n342 n330 U400/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M764 U400/a_25_64# n330 n342 VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M765 n342 n329 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M766 GND n350 n342 GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M767 n342 n330 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M768 VDD n266 U401/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M769 U401/a_18_54# U401/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M770 N395 n266 U401/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M771 U401/a_35_54# U401/a_2_6# N395 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M772 VDD G12 U401/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M773 U401/a_13_43# G12 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M774 GND n266 U401/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M775 U401/a_18_6# U401/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M776 N395 U401/a_2_6# U401/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M777 U401/a_35_6# n266 N395 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M778 GND G12 U401/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M779 U401/a_13_43# G12 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M780 VDD n259 U402/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M781 U402/a_18_54# U402/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M782 N394 n259 U402/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M783 U402/a_35_54# U402/a_2_6# N394 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M784 VDD G11 U402/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M785 U402/a_13_43# G11 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M786 GND n259 U402/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M787 U402/a_18_6# U402/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M788 N394 U402/a_2_6# U402/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M789 U402/a_35_6# n259 N394 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M790 GND G11 U402/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M791 U402/a_13_43# G11 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M792 VDD n241 U403/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M793 U403/a_18_54# U403/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M794 N393 U403/a_2_6# U403/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M795 U403/a_35_54# n241 N393 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M796 VDD n347 U403/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M797 U403/a_12_41# n347 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M798 GND n241 U403/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M799 U403/a_18_6# U403/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M800 N393 n241 U403/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M801 U403/a_35_6# U403/a_2_6# N393 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M802 GND n347 U403/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M803 U403/a_12_41# n347 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M804 VDD n252 U404/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M805 U404/a_18_54# U404/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M806 N392 n252 U404/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M807 U404/a_35_54# U404/a_2_6# N392 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M808 VDD G9 U404/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M809 U404/a_13_43# G9 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M810 GND n252 U404/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M811 U404/a_18_6# U404/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M812 N392 U404/a_2_6# U404/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M813 U404/a_35_6# n252 N392 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M814 GND G9 U404/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M815 U404/a_13_43# G9 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M816 n344 n227 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M817 n344 n227 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M818 n349 n327 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M819 VDD n239 n349 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M820 n349 n236 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M821 U406/a_9_6# n327 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M822 U406/a_14_6# n239 U406/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M823 n349 n236 U406/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M824 VDD n258 U407/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M825 U407/a_18_54# U407/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M826 N391 n258 U407/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M827 U407/a_35_54# U407/a_2_6# N391 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M828 VDD G8 U407/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M829 U407/a_13_43# G8 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M830 GND n258 U407/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M831 U407/a_18_6# U407/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M832 N391 U407/a_2_6# U407/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M833 U407/a_35_6# n258 N391 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M834 GND G8 U407/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M835 U407/a_13_43# G8 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M836 VDD n265 U408/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M837 U408/a_18_54# U408/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M838 N390 n265 U408/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M839 U408/a_35_54# U408/a_2_6# N390 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M840 VDD G7 U408/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M841 U408/a_13_43# G7 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M842 GND n265 U408/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M843 U408/a_18_6# U408/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M844 N390 U408/a_2_6# U408/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M845 U408/a_35_6# n265 N390 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M846 GND G7 U408/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M847 U408/a_13_43# G7 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M848 VDD n251 U409/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M849 U409/a_18_54# U409/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M850 N389 n251 U409/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M851 U409/a_35_54# U409/a_2_6# N389 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M852 VDD G6 U409/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M853 U409/a_13_43# G6 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M854 GND n251 U409/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M855 U409/a_18_6# U409/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M856 N389 U409/a_2_6# U409/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M857 U409/a_35_6# n251 N389 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M858 GND G6 U409/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M859 U409/a_13_43# G6 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M860 VDD n240 U410/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M861 U410/a_18_54# U410/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M862 N388 U410/a_2_6# U410/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M863 U410/a_35_54# n240 N388 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M864 VDD n357 U410/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M865 U410/a_12_41# n357 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M866 GND n240 U410/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M867 U410/a_18_6# U410/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M868 N388 n240 U410/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M869 U410/a_35_6# U410/a_2_6# N388 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M870 GND n357 U410/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M871 U410/a_12_41# n357 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M872 n353 n228 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M873 n353 n228 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M874 n358 n330 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M875 VDD n239 n358 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M876 n358 n237 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M877 U412/a_9_6# n330 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M878 U412/a_14_6# n239 U412/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M879 n358 n237 U412/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M880 VDD n250 U413/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M881 U413/a_18_54# U413/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M882 N387 n250 U413/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M883 U413/a_35_54# U413/a_2_6# N387 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M884 VDD G4 U413/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M885 U413/a_13_43# G4 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M886 GND n250 U413/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M887 U413/a_18_6# U413/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M888 N387 U413/a_2_6# U413/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M889 U413/a_35_6# n250 N387 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M890 GND G4 U413/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M891 U413/a_13_43# G4 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M892 VDD n246 U414/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M893 U414/a_18_54# U414/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M894 N386 n246 U414/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M895 U414/a_35_54# U414/a_2_6# N386 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M896 VDD G3 U414/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M897 U414/a_13_43# G3 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M898 GND n246 U414/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M899 U414/a_18_6# U414/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M900 N386 U414/a_2_6# U414/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M901 U414/a_35_6# n246 N386 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M902 GND G3 U414/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M903 U414/a_13_43# G3 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M904 VDD n278 U415/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M905 U415/a_18_54# U415/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M906 N385 n278 U415/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M907 U415/a_35_54# U415/a_2_6# N385 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M908 VDD G2 U415/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M909 U415/a_13_43# G2 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M910 GND n278 U415/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M911 U415/a_18_6# U415/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M912 N385 U415/a_2_6# U415/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M913 U415/a_35_6# n278 N385 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M914 GND G2 U415/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M915 U415/a_13_43# G2 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M916 VDD n272 U416/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M917 U416/a_18_54# U416/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M918 N384 n272 U416/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M919 U416/a_35_54# U416/a_2_6# N384 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M920 VDD G1 U416/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M921 U416/a_13_43# G1 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M922 GND n272 U416/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M923 U416/a_18_6# U416/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M924 N384 U416/a_2_6# U416/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M925 U416/a_35_6# n272 N384 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M926 GND G1 U416/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M927 U416/a_13_43# G1 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M928 n361 n229 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M929 n361 n229 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M930 n365 n330 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M931 VDD n329 n365 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M932 n365 n366 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M933 U418/a_9_6# n330 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M934 U418/a_14_6# n329 U418/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M935 n365 n366 U418/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M936 VDD n327 U419/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M937 U419/a_2_64# n327 VDD VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M938 U419/a_25_64# n350 U419/a_2_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M939 U419/a_2_64# n350 U419/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M940 n366 n332 U419/a_25_64# VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M941 U419/a_25_64# n332 n366 VDD pmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M942 n366 n327 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M943 GND n350 n366 GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M944 n366 n332 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M945 n332 n288 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M946 n332 n288 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M947 VDD n367 U421/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M948 U421/a_18_54# U421/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M949 n288 U421/a_2_6# U421/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M950 U421/a_35_54# n367 n288 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M951 VDD n368 U421/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M952 U421/a_12_41# n368 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M953 GND n367 U421/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M954 U421/a_18_6# U421/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M955 n288 n367 U421/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M956 U421/a_35_6# U421/a_2_6# n288 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M957 GND n368 U421/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M958 U421/a_12_41# n368 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M959 VDD n369 U422/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M960 U422/a_18_54# U422/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M961 n368 n369 U422/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M962 U422/a_35_54# U422/a_2_6# n368 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M963 VDD n370 U422/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M964 U422/a_13_43# n370 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M965 GND n369 U422/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M966 U422/a_18_6# U422/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M967 n368 U422/a_2_6# U422/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M968 U422/a_35_6# n369 n368 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M969 GND n370 U422/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M970 U422/a_13_43# n370 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M971 VDD G23 U423/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M972 U423/a_18_54# U423/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M973 n370 G23 U423/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M974 U423/a_35_54# U423/a_2_6# n370 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M975 VDD G19 U423/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M976 U423/a_13_43# G19 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M977 GND G23 U423/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M978 U423/a_18_6# U423/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M979 n370 U423/a_2_6# U423/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M980 U423/a_35_6# G23 n370 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M981 GND G19 U423/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M982 U423/a_13_43# G19 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M983 VDD G31 U424/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M984 U424/a_18_54# U424/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M985 n369 G31 U424/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M986 U424/a_35_54# U424/a_2_6# n369 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M987 VDD G27 U424/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M988 U424/a_13_43# G27 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M989 GND G31 U424/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M990 U424/a_18_6# U424/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M991 n369 U424/a_2_6# U424/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M992 U424/a_35_6# G31 n369 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M993 GND G27 U424/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M994 U424/a_13_43# G27 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M995 VDD n371 U425/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M996 U425/a_18_54# U425/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M997 n367 n371 U425/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M998 U425/a_35_54# U425/a_2_6# n367 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M999 VDD n372 U425/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1000 U425/a_13_43# n372 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1001 GND n371 U425/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1002 U425/a_18_6# U425/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1003 n367 U425/a_2_6# U425/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1004 U425/a_35_6# n371 n367 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1005 GND n372 U425/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1006 U425/a_13_43# n372 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1007 VDD n248 U426/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1008 U426/a_18_54# U426/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1009 n371 n248 U426/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1010 U426/a_35_54# U426/a_2_6# n371 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1011 VDD n374 U426/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1012 U426/a_13_43# n374 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1013 GND n248 U426/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1014 U426/a_18_6# U426/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1015 n371 U426/a_2_6# U426/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1016 U426/a_35_6# n248 n371 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1017 GND n374 U426/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1018 U426/a_13_43# n374 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1019 n376 n295 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1020 VDD n276 n376 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1021 n376 n298 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1022 U427/a_9_6# n295 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1023 U427/a_14_6# n276 U427/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1024 n376 n298 U427/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1025 n298 n307 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1026 n298 n307 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1027 n295 n340 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1028 n295 n340 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1029 n375 n294 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1030 VDD n282 n375 VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1031 n375 n297 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1032 U430/a_9_6# n294 GND GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1033 U430/a_14_6# n282 U430/a_9_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1034 n375 n297 U430/a_14_6# GND nmos W=0.75u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1035 n297 n316 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1036 n297 n316 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1037 VDD n377 U432/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1038 U432/a_18_54# U432/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1039 n316 U432/a_2_6# U432/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1040 U432/a_35_54# n377 n316 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1041 VDD n378 U432/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1042 U432/a_12_41# n378 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1043 GND n377 U432/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1044 U432/a_18_6# U432/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1045 n316 n377 U432/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1046 U432/a_35_6# U432/a_2_6# n316 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1047 GND n378 U432/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1048 U432/a_12_41# n378 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1049 VDD n379 U433/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1050 U433/a_18_54# U433/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1051 n378 n379 U433/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1052 U433/a_35_54# U433/a_2_6# n378 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1053 VDD n380 U433/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1054 U433/a_13_43# n380 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1055 GND n379 U433/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1056 U433/a_18_6# U433/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1057 n378 U433/a_2_6# U433/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1058 U433/a_35_6# n379 n378 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1059 GND n380 U433/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1060 U433/a_13_43# n380 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1061 VDD G14 U434/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1062 U434/a_18_54# U434/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1063 n380 U434/a_2_6# U434/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1064 U434/a_35_54# G14 n380 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1065 VDD n347 U434/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1066 U434/a_12_41# n347 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1067 GND G14 U434/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1068 U434/a_18_6# U434/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1069 n380 G14 U434/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1070 U434/a_35_6# U434/a_2_6# n380 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1071 GND n347 U434/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1072 U434/a_12_41# n347 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1073 n347 G10 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1074 n347 G10 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1075 VDD G6 U436/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1076 U436/a_18_54# U436/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1077 n379 G6 U436/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1078 U436/a_35_54# U436/a_2_6# n379 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1079 VDD G2 U436/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1080 U436/a_13_43# G2 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1081 GND G6 U436/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1082 U436/a_18_6# U436/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1083 n379 U436/a_2_6# U436/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1084 U436/a_35_6# G6 n379 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1085 GND G2 U436/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1086 U436/a_13_43# G2 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1087 VDD n381 U437/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1088 U437/a_18_54# U437/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1089 n377 n381 U437/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1090 U437/a_35_54# U437/a_2_6# n377 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1091 VDD n382 U437/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1092 U437/a_13_43# n382 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1093 GND n381 U437/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1094 U437/a_18_6# U437/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1095 n377 U437/a_2_6# U437/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1096 U437/a_35_6# n381 n377 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1097 GND n382 U437/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1098 U437/a_13_43# n382 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1099 VDD n257 U438/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1100 U438/a_18_54# U438/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1101 n381 n257 U438/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1102 U438/a_35_54# U438/a_2_6# n381 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1103 VDD n384 U438/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1104 U438/a_13_43# n384 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1105 GND n257 U438/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1106 U438/a_18_6# U438/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1107 n381 U438/a_2_6# U438/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1108 U438/a_35_6# n257 n381 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1109 GND n384 U438/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1110 U438/a_13_43# n384 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1111 VDD n385 U439/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1112 U439/a_18_54# U439/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1113 n307 U439/a_2_6# U439/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1114 U439/a_35_54# n385 n307 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1115 VDD n386 U439/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1116 U439/a_12_41# n386 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1117 GND n385 U439/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1118 U439/a_18_6# U439/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1119 n307 n385 U439/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1120 U439/a_35_6# U439/a_2_6# n307 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1121 GND n386 U439/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1122 U439/a_12_41# n386 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1123 VDD n387 U440/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1124 U440/a_18_54# U440/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1125 n386 n387 U440/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1126 U440/a_35_54# U440/a_2_6# n386 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1127 VDD n388 U440/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1128 U440/a_13_43# n388 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1129 GND n387 U440/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1130 U440/a_18_6# U440/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1131 n386 U440/a_2_6# U440/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1132 U440/a_35_6# n387 n386 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1133 GND n388 U440/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1134 U440/a_13_43# n388 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1135 VDD G16 U441/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1136 U441/a_18_54# U441/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1137 n388 G16 U441/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1138 U441/a_35_54# U441/a_2_6# n388 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1139 VDD G12 U441/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1140 U441/a_13_43# G12 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1141 GND G16 U441/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1142 U441/a_18_6# U441/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1143 n388 U441/a_2_6# U441/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1144 U441/a_35_6# G16 n388 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1145 GND G12 U441/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1146 U441/a_13_43# G12 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1147 VDD G8 U442/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1148 U442/a_18_54# U442/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1149 n387 G8 U442/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1150 U442/a_35_54# U442/a_2_6# n387 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1151 VDD G4 U442/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1152 U442/a_13_43# G4 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1153 GND G8 U442/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1154 U442/a_18_6# U442/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1155 n387 U442/a_2_6# U442/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1156 U442/a_35_6# G8 n387 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1157 GND G4 U442/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1158 U442/a_13_43# G4 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1159 VDD n389 U443/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1160 U443/a_18_54# U443/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1161 n385 n389 U443/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1162 U443/a_35_54# U443/a_2_6# n385 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1163 VDD n390 U443/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1164 U443/a_13_43# n390 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1165 GND n389 U443/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1166 U443/a_18_6# U443/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1167 n385 U443/a_2_6# U443/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1168 U443/a_35_6# n389 n385 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1169 GND n390 U443/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1170 U443/a_13_43# n390 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1171 VDD n242 U444/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1172 U444/a_18_54# U444/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1173 n389 n242 U444/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1174 U444/a_35_54# U444/a_2_6# n389 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1175 VDD n384 U444/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1176 U444/a_13_43# n384 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1177 GND n242 U444/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1178 U444/a_18_6# U444/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1179 n389 U444/a_2_6# U444/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1180 U444/a_35_6# n242 n389 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1181 GND n384 U444/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1182 U444/a_13_43# n384 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1183 VDD n392 U445/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1184 U445/a_18_54# U445/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1185 n384 U445/a_2_6# U445/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1186 U445/a_35_54# n392 n384 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1187 VDD n393 U445/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1188 U445/a_12_41# n393 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1189 GND n392 U445/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1190 U445/a_18_6# U445/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1191 n384 n392 U445/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1192 U445/a_35_6# U445/a_2_6# n384 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1193 GND n393 U445/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1194 U445/a_12_41# n393 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1195 VDD G32 U446/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1196 U446/a_18_54# U446/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1197 n393 G32 U446/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1198 U446/a_35_54# U446/a_2_6# n393 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1199 VDD G31 U446/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1200 U446/a_13_43# G31 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1201 GND G32 U446/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1202 U446/a_18_6# U446/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1203 n393 U446/a_2_6# U446/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1204 U446/a_35_6# G32 n393 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1205 GND G31 U446/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1206 U446/a_13_43# G31 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1207 VDD G29 U447/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1208 U447/a_18_54# U447/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1209 n392 U447/a_2_6# U447/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1210 U447/a_35_54# G29 n392 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1211 VDD G30 U447/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1212 U447/a_12_41# G30 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1213 GND G29 U447/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1214 U447/a_18_6# U447/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1215 n392 G29 U447/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1216 U447/a_35_6# U447/a_2_6# n392 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1217 GND G30 U447/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1218 U447/a_12_41# G30 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1219 VDD n394 U448/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1220 U448/a_18_54# U448/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1221 n340 U448/a_2_6# U448/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1222 U448/a_35_54# n394 n340 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1223 VDD n395 U448/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1224 U448/a_12_41# n395 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1225 GND n394 U448/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1226 U448/a_18_6# U448/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1227 n340 n394 U448/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1228 U448/a_35_6# U448/a_2_6# n340 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1229 GND n395 U448/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1230 U448/a_12_41# n395 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1231 VDD n396 U449/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1232 U449/a_18_54# U449/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1233 n395 n396 U449/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1234 U449/a_35_54# U449/a_2_6# n395 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1235 VDD n397 U449/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1236 U449/a_13_43# n397 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1237 GND n396 U449/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1238 U449/a_18_6# U449/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1239 n395 U449/a_2_6# U449/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1240 U449/a_35_6# n396 n395 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1241 GND n397 U449/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1242 U449/a_13_43# n397 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1243 VDD n339 U450/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1244 U450/a_18_54# U450/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1245 n397 U450/a_2_6# U450/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1246 U450/a_35_54# n339 n397 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1247 VDD G1 U450/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1248 U450/a_12_41# G1 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1249 GND n339 U450/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1250 U450/a_18_6# U450/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1251 n397 n339 U450/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1252 U450/a_35_6# U450/a_2_6# n397 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1253 GND G1 U450/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1254 U450/a_12_41# G1 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1255 n339 G13 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1256 n339 G13 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1257 VDD G9 U452/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1258 U452/a_18_54# U452/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1259 n396 U452/a_2_6# U452/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1260 U452/a_35_54# G9 n396 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1261 VDD n357 U452/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1262 U452/a_12_41# n357 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1263 GND G9 U452/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1264 U452/a_18_6# U452/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1265 n396 G9 U452/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1266 U452/a_35_6# U452/a_2_6# n396 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1267 GND n357 U452/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1268 U452/a_12_41# n357 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1269 n357 G5 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1270 n357 G5 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1271 VDD n398 U454/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1272 U454/a_18_54# U454/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1273 n394 n398 U454/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1274 U454/a_35_54# U454/a_2_6# n394 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1275 VDD n399 U454/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1276 U454/a_13_43# n399 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1277 GND n398 U454/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1278 U454/a_18_6# U454/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1279 n394 U454/a_2_6# U454/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1280 U454/a_35_6# n398 n394 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1281 GND n399 U454/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1282 U454/a_13_43# n399 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1283 VDD n264 U455/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1284 U455/a_18_54# U455/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1285 n398 n264 U455/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1286 U455/a_35_54# U455/a_2_6# n398 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1287 VDD n390 U455/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1288 U455/a_13_43# n390 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1289 GND n264 U455/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1290 U455/a_18_6# U455/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1291 n398 U455/a_2_6# U455/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1292 U455/a_35_6# n264 n398 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1293 GND n390 U455/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1294 U455/a_13_43# n390 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1295 VDD n401 U456/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1296 U456/a_18_54# U456/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1297 n390 U456/a_2_6# U456/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1298 U456/a_35_54# n401 n390 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1299 VDD n402 U456/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1300 U456/a_12_41# n402 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1301 GND n401 U456/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1302 U456/a_18_6# U456/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1303 n390 n401 U456/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1304 U456/a_35_6# U456/a_2_6# n390 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1305 GND n402 U456/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1306 U456/a_12_41# n402 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1307 VDD G24 U457/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1308 U457/a_18_54# U457/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1309 n402 G24 U457/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1310 U457/a_35_54# U457/a_2_6# n402 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1311 VDD G23 U457/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1312 U457/a_13_43# G23 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1313 GND G24 U457/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1314 U457/a_18_6# U457/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1315 n402 U457/a_2_6# U457/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1316 U457/a_35_6# G24 n402 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1317 GND G23 U457/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1318 U457/a_13_43# G23 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1319 VDD G21 U458/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1320 U458/a_18_54# U458/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1321 n401 U458/a_2_6# U458/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1322 U458/a_35_54# G21 n401 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1323 VDD G22 U458/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1324 U458/a_12_41# G22 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1325 GND G21 U458/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1326 U458/a_18_6# U458/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1327 n401 G21 U458/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1328 U458/a_35_6# U458/a_2_6# n401 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1329 GND G22 U458/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1330 U458/a_12_41# G22 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1331 n294 n336 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1332 n294 n336 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1333 VDD n403 U460/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1334 U460/a_18_54# U460/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1335 n336 U460/a_2_6# U460/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1336 U460/a_35_54# n403 n336 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1337 VDD n404 U460/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1338 U460/a_12_41# n404 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1339 GND n403 U460/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1340 U460/a_18_6# U460/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1341 n336 n403 U460/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1342 U460/a_35_6# U460/a_2_6# n336 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1343 GND n404 U460/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1344 U460/a_12_41# n404 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1345 VDD n405 U461/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1346 U461/a_18_54# U461/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1347 n404 n405 U461/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1348 U461/a_35_54# U461/a_2_6# n404 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1349 VDD n406 U461/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1350 U461/a_13_43# n406 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1351 GND n405 U461/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1352 U461/a_18_6# U461/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1353 n404 U461/a_2_6# U461/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1354 U461/a_35_6# n405 n404 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1355 GND n406 U461/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1356 U461/a_13_43# n406 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1357 VDD G15 U462/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1358 U462/a_18_54# U462/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1359 n406 G15 U462/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1360 U462/a_35_54# U462/a_2_6# n406 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1361 VDD G11 U462/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1362 U462/a_13_43# G11 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1363 GND G15 U462/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1364 U462/a_18_6# U462/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1365 n406 U462/a_2_6# U462/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1366 U462/a_35_6# G15 n406 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1367 GND G11 U462/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1368 U462/a_13_43# G11 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1369 VDD G7 U463/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1370 U463/a_18_54# U463/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1371 n405 G7 U463/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1372 U463/a_35_54# U463/a_2_6# n405 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1373 VDD G3 U463/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1374 U463/a_13_43# G3 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1375 GND G7 U463/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1376 U463/a_18_6# U463/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1377 n405 U463/a_2_6# U463/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1378 U463/a_35_6# G7 n405 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1379 GND G3 U463/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1380 U463/a_13_43# G3 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1381 VDD n407 U464/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1382 U464/a_18_54# U464/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1383 n403 n407 U464/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1384 U464/a_35_54# U464/a_2_6# n403 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1385 VDD n399 U464/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1386 U464/a_13_43# n399 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1387 GND n407 U464/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1388 U464/a_18_6# U464/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1389 n403 U464/a_2_6# U464/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1390 U464/a_35_6# n407 n403 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1391 GND n399 U464/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1392 U464/a_13_43# n399 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1393 VDD n408 U465/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1394 U465/a_18_54# U465/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1395 n399 U465/a_2_6# U465/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1396 U465/a_35_54# n408 n399 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1397 VDD n409 U465/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1398 U465/a_12_41# n409 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1399 GND n408 U465/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1400 U465/a_18_6# U465/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1401 n399 n408 U465/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1402 U465/a_35_6# U465/a_2_6# n399 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1403 GND n409 U465/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1404 U465/a_12_41# n409 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1405 VDD G20 U466/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1406 U466/a_18_54# U466/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1407 n409 G20 U466/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1408 U466/a_35_54# U466/a_2_6# n409 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1409 VDD G19 U466/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1410 U466/a_13_43# G19 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1411 GND G20 U466/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1412 U466/a_18_6# U466/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1413 n409 U466/a_2_6# U466/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1414 U466/a_35_6# G20 n409 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1415 GND G19 U466/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1416 U466/a_13_43# G19 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1417 VDD G17 U467/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1418 U467/a_18_54# U467/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1419 n408 U467/a_2_6# U467/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1420 U467/a_35_54# G17 n408 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1421 VDD G18 U467/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1422 U467/a_12_41# G18 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1423 GND G17 U467/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1424 U467/a_18_6# U467/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1425 n408 G17 U467/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1426 U467/a_35_6# U467/a_2_6# n408 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1427 GND G18 U467/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1428 U467/a_12_41# G18 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1429 VDD n249 U468/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1430 U468/a_18_54# U468/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1431 n407 n249 U468/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1432 U468/a_35_54# U468/a_2_6# n407 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1433 VDD n382 U468/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1434 U468/a_13_43# n382 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1435 GND n249 U468/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1436 U468/a_18_6# U468/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1437 n407 U468/a_2_6# U468/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1438 U468/a_35_6# n249 n407 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1439 GND n382 U468/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1440 U468/a_13_43# n382 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1441 VDD n411 U469/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1442 U469/a_18_54# U469/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1443 n382 U469/a_2_6# U469/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1444 U469/a_35_54# n411 n382 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1445 VDD n412 U469/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1446 U469/a_12_41# n412 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1447 GND n411 U469/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1448 U469/a_18_6# U469/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1449 n382 n411 U469/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1450 U469/a_35_6# U469/a_2_6# n382 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1451 GND n412 U469/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1452 U469/a_12_41# n412 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1453 VDD G28 U470/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1454 U470/a_18_54# U470/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1455 n412 G28 U470/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1456 U470/a_35_54# U470/a_2_6# n412 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1457 VDD G27 U470/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1458 U470/a_13_43# G27 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1459 GND G28 U470/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1460 U470/a_18_6# U470/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1461 n412 U470/a_2_6# U470/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1462 U470/a_35_6# G28 n412 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1463 GND G27 U470/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1464 U470/a_13_43# G27 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1465 VDD G25 U471/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1466 U471/a_18_54# U471/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1467 n411 U471/a_2_6# U471/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1468 U471/a_35_54# G25 n411 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1469 VDD G26 U471/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1470 U471/a_12_41# G26 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1471 GND G25 U471/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1472 U471/a_18_6# U471/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1473 n411 G25 U471/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1474 U471/a_35_6# U471/a_2_6# n411 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1475 GND G26 U471/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1476 U471/a_12_41# G26 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1477 n327 n292 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1478 n327 n292 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1479 VDD n413 U473/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1480 U473/a_18_54# U473/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1481 n292 U473/a_2_6# U473/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1482 U473/a_35_54# n413 n292 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1483 VDD n414 U473/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1484 U473/a_12_41# n414 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1485 GND n413 U473/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1486 U473/a_18_6# U473/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1487 n292 n413 U473/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1488 U473/a_35_6# U473/a_2_6# n292 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1489 GND n414 U473/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1490 U473/a_12_41# n414 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1491 VDD n415 U474/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1492 U474/a_18_54# U474/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1493 n414 n415 U474/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1494 U474/a_35_54# U474/a_2_6# n414 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1495 VDD n416 U474/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1496 U474/a_13_43# n416 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1497 GND n415 U474/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1498 U474/a_18_6# U474/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1499 n414 U474/a_2_6# U474/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1500 U474/a_35_6# n415 n414 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1501 GND n416 U474/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1502 U474/a_13_43# n416 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1503 VDD G21 U475/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1504 U475/a_18_54# U475/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1505 n416 G21 U475/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1506 U475/a_35_54# U475/a_2_6# n416 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1507 VDD G17 U475/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1508 U475/a_13_43# G17 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1509 GND G21 U475/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1510 U475/a_18_6# U475/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1511 n416 U475/a_2_6# U475/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1512 U475/a_35_6# G21 n416 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1513 GND G17 U475/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1514 U475/a_13_43# G17 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1515 VDD G29 U476/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1516 U476/a_18_54# U476/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1517 n415 G29 U476/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1518 U476/a_35_54# U476/a_2_6# n415 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1519 VDD G25 U476/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1520 U476/a_13_43# G25 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1521 GND G29 U476/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1522 U476/a_18_6# U476/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1523 n415 U476/a_2_6# U476/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1524 U476/a_35_6# G29 n415 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1525 GND G25 U476/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1526 U476/a_13_43# G25 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1527 VDD n417 U477/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1528 U477/a_18_54# U477/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1529 n413 n417 U477/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1530 U477/a_35_54# U477/a_2_6# n413 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1531 VDD n372 U477/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1532 U477/a_13_43# n372 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1533 GND n417 U477/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1534 U477/a_18_6# U477/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1535 n413 U477/a_2_6# U477/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1536 U477/a_35_6# n417 n413 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1537 GND n372 U477/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1538 U477/a_13_43# n372 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1539 VDD n418 U478/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1540 U478/a_18_54# U478/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1541 n372 U478/a_2_6# U478/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1542 U478/a_35_54# n418 n372 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1543 VDD n419 U478/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1544 U478/a_12_41# n419 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1545 GND n418 U478/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1546 U478/a_18_6# U478/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1547 n372 n418 U478/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1548 U478/a_35_6# U478/a_2_6# n372 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1549 GND n419 U478/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1550 U478/a_12_41# n419 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1551 VDD G4 U479/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1552 U479/a_18_54# U479/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1553 n419 G4 U479/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1554 U479/a_35_54# U479/a_2_6# n419 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1555 VDD G3 U479/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1556 U479/a_13_43# G3 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1557 GND G4 U479/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1558 U479/a_18_6# U479/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1559 n419 U479/a_2_6# U479/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1560 U479/a_35_6# G4 n419 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1561 GND G3 U479/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1562 U479/a_13_43# G3 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1563 VDD G1 U480/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1564 U480/a_18_54# U480/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1565 n418 U480/a_2_6# U480/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1566 U480/a_35_54# G1 n418 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1567 VDD G2 U480/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1568 U480/a_12_41# G2 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1569 GND G1 U480/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1570 U480/a_18_6# U480/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1571 n418 G1 U480/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1572 U480/a_35_6# U480/a_2_6# n418 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1573 GND G2 U480/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1574 U480/a_12_41# G2 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1575 VDD n244 U481/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1576 U481/a_18_54# U481/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1577 n417 n244 U481/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1578 U481/a_35_54# U481/a_2_6# n417 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1579 VDD n421 U481/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1580 U481/a_13_43# n421 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1581 GND n244 U481/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1582 U481/a_18_6# U481/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1583 n417 U481/a_2_6# U481/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1584 U481/a_35_6# n244 n417 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1585 GND n421 U481/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1586 U481/a_13_43# n421 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1587 n329 n286 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1588 n329 n286 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1589 VDD n422 U483/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1590 U483/a_18_54# U483/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1591 n286 U483/a_2_6# U483/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1592 U483/a_35_54# n422 n286 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1593 VDD n423 U483/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1594 U483/a_12_41# n423 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1595 GND n422 U483/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1596 U483/a_18_6# U483/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1597 n286 n422 U483/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1598 U483/a_35_6# U483/a_2_6# n286 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1599 GND n423 U483/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1600 U483/a_12_41# n423 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1601 VDD n424 U484/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1602 U484/a_18_54# U484/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1603 n423 n424 U484/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1604 U484/a_35_54# U484/a_2_6# n423 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1605 VDD n425 U484/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1606 U484/a_13_43# n425 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1607 GND n424 U484/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1608 U484/a_18_6# U484/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1609 n423 U484/a_2_6# U484/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1610 U484/a_35_6# n424 n423 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1611 GND n425 U484/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1612 U484/a_13_43# n425 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1613 VDD G24 U485/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1614 U485/a_18_54# U485/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1615 n425 G24 U485/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1616 U485/a_35_54# U485/a_2_6# n425 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1617 VDD G20 U485/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1618 U485/a_13_43# G20 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1619 GND G24 U485/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1620 U485/a_18_6# U485/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1621 n425 U485/a_2_6# U485/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1622 U485/a_35_6# G24 n425 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1623 GND G20 U485/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1624 U485/a_13_43# G20 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1625 VDD G32 U486/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1626 U486/a_18_54# U486/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1627 n424 G32 U486/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1628 U486/a_35_54# U486/a_2_6# n424 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1629 VDD G28 U486/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1630 U486/a_13_43# G28 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1631 GND G32 U486/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1632 U486/a_18_6# U486/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1633 n424 U486/a_2_6# U486/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1634 U486/a_35_6# G32 n424 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1635 GND G28 U486/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1636 U486/a_13_43# G28 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1637 VDD n426 U487/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1638 U487/a_18_54# U487/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1639 n422 n426 U487/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1640 U487/a_35_54# U487/a_2_6# n422 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1641 VDD n421 U487/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1642 U487/a_13_43# n421 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1643 GND n426 U487/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1644 U487/a_18_6# U487/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1645 n422 U487/a_2_6# U487/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1646 U487/a_35_6# n426 n422 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1647 GND n421 U487/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1648 U487/a_13_43# n421 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1649 VDD n427 U488/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1650 U488/a_18_54# U488/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1651 n421 U488/a_2_6# U488/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1652 U488/a_35_54# n427 n421 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1653 VDD n428 U488/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1654 U488/a_12_41# n428 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1655 GND n427 U488/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1656 U488/a_18_6# U488/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1657 n421 n427 U488/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1658 U488/a_35_6# U488/a_2_6# n421 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1659 GND n428 U488/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1660 U488/a_12_41# n428 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1661 VDD G8 U489/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1662 U489/a_18_54# U489/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1663 n428 G8 U489/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1664 U489/a_35_54# U489/a_2_6# n428 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1665 VDD G7 U489/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1666 U489/a_13_43# G7 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1667 GND G8 U489/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1668 U489/a_18_6# U489/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1669 n428 U489/a_2_6# U489/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1670 U489/a_35_6# G8 n428 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1671 GND G7 U489/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1672 U489/a_13_43# G7 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1673 VDD G5 U490/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1674 U490/a_18_54# U490/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1675 n427 U490/a_2_6# U490/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1676 U490/a_35_54# G5 n427 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1677 VDD G6 U490/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1678 U490/a_12_41# G6 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1679 GND G5 U490/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1680 U490/a_18_6# U490/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1681 n427 G5 U490/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1682 U490/a_35_6# U490/a_2_6# n427 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1683 GND G6 U490/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1684 U490/a_12_41# G6 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1685 VDD n245 U491/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1686 U491/a_18_54# U491/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1687 n426 n245 U491/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1688 U491/a_35_54# U491/a_2_6# n426 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1689 VDD n430 U491/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1690 U491/a_13_43# n430 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1691 GND n245 U491/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1692 U491/a_18_6# U491/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1693 n426 U491/a_2_6# U491/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1694 U491/a_35_6# n245 n426 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1695 GND n430 U491/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1696 U491/a_13_43# n430 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1697 n330 n290 VDD VDD pmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1698 n330 n290 GND GND nmos W=0.25u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1699 VDD n431 U493/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1700 U493/a_18_54# U493/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1701 n290 U493/a_2_6# U493/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1702 U493/a_35_54# n431 n290 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1703 VDD n432 U493/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1704 U493/a_12_41# n432 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1705 GND n431 U493/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1706 U493/a_18_6# U493/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1707 n290 n431 U493/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1708 U493/a_35_6# U493/a_2_6# n290 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1709 GND n432 U493/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1710 U493/a_12_41# n432 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1711 VDD n433 U494/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1712 U494/a_18_54# U494/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1713 n432 n433 U494/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1714 U494/a_35_54# U494/a_2_6# n432 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1715 VDD n434 U494/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1716 U494/a_13_43# n434 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1717 GND n433 U494/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1718 U494/a_18_6# U494/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1719 n432 U494/a_2_6# U494/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1720 U494/a_35_6# n433 n432 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1721 GND n434 U494/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1722 U494/a_13_43# n434 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1723 VDD G22 U495/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1724 U495/a_18_54# U495/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1725 n434 G22 U495/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1726 U495/a_35_54# U495/a_2_6# n434 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1727 VDD G18 U495/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1728 U495/a_13_43# G18 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1729 GND G22 U495/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1730 U495/a_18_6# U495/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1731 n434 U495/a_2_6# U495/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1732 U495/a_35_6# G22 n434 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1733 GND G18 U495/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1734 U495/a_13_43# G18 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1735 VDD G30 U496/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1736 U496/a_18_54# U496/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1737 n433 G30 U496/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1738 U496/a_35_54# U496/a_2_6# n433 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1739 VDD G26 U496/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1740 U496/a_13_43# G26 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1741 GND G30 U496/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1742 U496/a_18_6# U496/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1743 n433 U496/a_2_6# U496/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1744 U496/a_35_6# G30 n433 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1745 GND G26 U496/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1746 U496/a_13_43# G26 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1747 VDD n435 U497/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1748 U497/a_18_54# U497/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1749 n431 n435 U497/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1750 U497/a_35_54# U497/a_2_6# n431 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1751 VDD n374 U497/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1752 U497/a_13_43# n374 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1753 GND n435 U497/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1754 U497/a_18_6# U497/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1755 n431 U497/a_2_6# U497/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1756 U497/a_35_6# n435 n431 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1757 GND n374 U497/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1758 U497/a_13_43# n374 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1759 VDD n436 U498/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1760 U498/a_18_54# U498/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1761 n374 U498/a_2_6# U498/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1762 U498/a_35_54# n436 n374 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1763 VDD n437 U498/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1764 U498/a_12_41# n437 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1765 GND n436 U498/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1766 U498/a_18_6# U498/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1767 n374 n436 U498/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1768 U498/a_35_6# U498/a_2_6# n374 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1769 GND n437 U498/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1770 U498/a_12_41# n437 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1771 VDD G9 U499/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1772 U499/a_18_54# U499/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1773 n437 G9 U499/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1774 U499/a_35_54# U499/a_2_6# n437 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1775 VDD G12 U499/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1776 U499/a_13_43# G12 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1777 GND G9 U499/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1778 U499/a_18_6# U499/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1779 n437 U499/a_2_6# U499/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1780 U499/a_35_6# G9 n437 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1781 GND G12 U499/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1782 U499/a_13_43# G12 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1783 VDD G10 U500/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1784 U500/a_18_54# U500/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1785 n436 U500/a_2_6# U500/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1786 U500/a_35_54# G10 n436 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1787 VDD G11 U500/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1788 U500/a_12_41# G11 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1789 GND G10 U500/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1790 U500/a_18_6# U500/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1791 n436 G10 U500/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1792 U500/a_35_6# U500/a_2_6# n436 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1793 GND G11 U500/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1794 U500/a_12_41# G11 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1795 VDD n243 U501/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1796 U501/a_18_54# U501/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1797 n435 n243 U501/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1798 U501/a_35_54# U501/a_2_6# n435 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1799 VDD n430 U501/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1800 U501/a_13_43# n430 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1801 GND n243 U501/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1802 U501/a_18_6# U501/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1803 n435 U501/a_2_6# U501/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1804 U501/a_35_6# n243 n435 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1805 GND n430 U501/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1806 U501/a_13_43# n430 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1807 VDD n439 U502/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1808 U502/a_18_54# U502/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1809 n430 U502/a_2_6# U502/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1810 U502/a_35_54# n439 n430 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1811 VDD n440 U502/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1812 U502/a_12_41# n440 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1813 GND n439 U502/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1814 U502/a_18_6# U502/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1815 n430 n439 U502/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1816 U502/a_35_6# U502/a_2_6# n430 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1817 GND n440 U502/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1818 U502/a_12_41# n440 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1819 VDD G16 U503/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1820 U503/a_18_54# U503/a_13_43# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1821 n440 G16 U503/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1822 U503/a_35_54# U503/a_2_6# n440 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1823 VDD G15 U503/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1824 U503/a_13_43# G15 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1825 GND G16 U503/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1826 U503/a_18_6# U503/a_13_43# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1827 n440 U503/a_2_6# U503/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1828 U503/a_35_6# G16 n440 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1829 GND G15 U503/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1830 U503/a_13_43# G15 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1831 VDD G13 U504/a_2_6# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1832 U504/a_18_54# U504/a_12_41# VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1833 n439 U504/a_2_6# U504/a_18_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1834 U504/a_35_54# G13 n439 VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1835 VDD G14 U504/a_35_54# VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1836 U504/a_12_41# G14 VDD VDD pmos W=1u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1837 GND G13 U504/a_2_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1838 U504/a_18_6# U504/a_12_41# GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1839 n439 G13 U504/a_18_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1840 U504/a_35_6# U504/a_2_6# n439 GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1841 GND G14 U504/a_35_6# GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
M1842 U504/a_12_41# G14 GND GND nmos W=0.5u L=0.05u AD=0p PD=0u AS=0p PS=0u 
.ENDS

